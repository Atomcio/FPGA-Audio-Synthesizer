library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package sine_lut_pkg is
  constant LUT_SIZE : integer := 4096;
  type sine_lut_t is array (0 to LUT_SIZE-1) of signed(15 downto 0);
  constant sine_lut : sine_lut_t := (
    0 => to_signed(0, 16),
    1 => to_signed(50, 16),
    2 => to_signed(100, 16),
    3 => to_signed(150, 16),
    4 => to_signed(201, 16),
    5 => to_signed(251, 16),
    6 => to_signed(301, 16),
    7 => to_signed(351, 16),
    8 => to_signed(402, 16),
    9 => to_signed(452, 16),
    10 => to_signed(502, 16),
    11 => to_signed(552, 16),
    12 => to_signed(603, 16),
    13 => to_signed(653, 16),
    14 => to_signed(703, 16),
    15 => to_signed(753, 16),
    16 => to_signed(804, 16),
    17 => to_signed(854, 16),
    18 => to_signed(904, 16),
    19 => to_signed(954, 16),
    20 => to_signed(1005, 16),
    21 => to_signed(1055, 16),
    22 => to_signed(1105, 16),
    23 => to_signed(1155, 16),
    24 => to_signed(1206, 16),
    25 => to_signed(1256, 16),
    26 => to_signed(1306, 16),
    27 => to_signed(1356, 16),
    28 => to_signed(1406, 16),
    29 => to_signed(1457, 16),
    30 => to_signed(1507, 16),
    31 => to_signed(1557, 16),
    32 => to_signed(1607, 16),
    33 => to_signed(1658, 16),
    34 => to_signed(1708, 16),
    35 => to_signed(1758, 16),
    36 => to_signed(1808, 16),
    37 => to_signed(1858, 16),
    38 => to_signed(1908, 16),
    39 => to_signed(1959, 16),
    40 => to_signed(2009, 16),
    41 => to_signed(2059, 16),
    42 => to_signed(2109, 16),
    43 => to_signed(2159, 16),
    44 => to_signed(2209, 16),
    45 => to_signed(2260, 16),
    46 => to_signed(2310, 16),
    47 => to_signed(2360, 16),
    48 => to_signed(2410, 16),
    49 => to_signed(2460, 16),
    50 => to_signed(2510, 16),
    51 => to_signed(2560, 16),
    52 => to_signed(2610, 16),
    53 => to_signed(2661, 16),
    54 => to_signed(2711, 16),
    55 => to_signed(2761, 16),
    56 => to_signed(2811, 16),
    57 => to_signed(2861, 16),
    58 => to_signed(2911, 16),
    59 => to_signed(2961, 16),
    60 => to_signed(3011, 16),
    61 => to_signed(3061, 16),
    62 => to_signed(3111, 16),
    63 => to_signed(3161, 16),
    64 => to_signed(3211, 16),
    65 => to_signed(3261, 16),
    66 => to_signed(3311, 16),
    67 => to_signed(3361, 16),
    68 => to_signed(3411, 16),
    69 => to_signed(3461, 16),
    70 => to_signed(3511, 16),
    71 => to_signed(3561, 16),
    72 => to_signed(3611, 16),
    73 => to_signed(3661, 16),
    74 => to_signed(3711, 16),
    75 => to_signed(3761, 16),
    76 => to_signed(3811, 16),
    77 => to_signed(3861, 16),
    78 => to_signed(3911, 16),
    79 => to_signed(3961, 16),
    80 => to_signed(4011, 16),
    81 => to_signed(4060, 16),
    82 => to_signed(4110, 16),
    83 => to_signed(4160, 16),
    84 => to_signed(4210, 16),
    85 => to_signed(4260, 16),
    86 => to_signed(4310, 16),
    87 => to_signed(4359, 16),
    88 => to_signed(4409, 16),
    89 => to_signed(4459, 16),
    90 => to_signed(4509, 16),
    91 => to_signed(4559, 16),
    92 => to_signed(4608, 16),
    93 => to_signed(4658, 16),
    94 => to_signed(4708, 16),
    95 => to_signed(4758, 16),
    96 => to_signed(4807, 16),
    97 => to_signed(4857, 16),
    98 => to_signed(4907, 16),
    99 => to_signed(4957, 16),
    100 => to_signed(5006, 16),
    101 => to_signed(5056, 16),
    102 => to_signed(5106, 16),
    103 => to_signed(5155, 16),
    104 => to_signed(5205, 16),
    105 => to_signed(5254, 16),
    106 => to_signed(5304, 16),
    107 => to_signed(5354, 16),
    108 => to_signed(5403, 16),
    109 => to_signed(5453, 16),
    110 => to_signed(5502, 16),
    111 => to_signed(5552, 16),
    112 => to_signed(5601, 16),
    113 => to_signed(5651, 16),
    114 => to_signed(5700, 16),
    115 => to_signed(5750, 16),
    116 => to_signed(5799, 16),
    117 => to_signed(5849, 16),
    118 => to_signed(5898, 16),
    119 => to_signed(5948, 16),
    120 => to_signed(5997, 16),
    121 => to_signed(6047, 16),
    122 => to_signed(6096, 16),
    123 => to_signed(6145, 16),
    124 => to_signed(6195, 16),
    125 => to_signed(6244, 16),
    126 => to_signed(6293, 16),
    127 => to_signed(6343, 16),
    128 => to_signed(6392, 16),
    129 => to_signed(6441, 16),
    130 => to_signed(6491, 16),
    131 => to_signed(6540, 16),
    132 => to_signed(6589, 16),
    133 => to_signed(6638, 16),
    134 => to_signed(6688, 16),
    135 => to_signed(6737, 16),
    136 => to_signed(6786, 16),
    137 => to_signed(6835, 16),
    138 => to_signed(6884, 16),
    139 => to_signed(6933, 16),
    140 => to_signed(6982, 16),
    141 => to_signed(7032, 16),
    142 => to_signed(7081, 16),
    143 => to_signed(7130, 16),
    144 => to_signed(7179, 16),
    145 => to_signed(7228, 16),
    146 => to_signed(7277, 16),
    147 => to_signed(7326, 16),
    148 => to_signed(7375, 16),
    149 => to_signed(7424, 16),
    150 => to_signed(7473, 16),
    151 => to_signed(7522, 16),
    152 => to_signed(7571, 16),
    153 => to_signed(7619, 16),
    154 => to_signed(7668, 16),
    155 => to_signed(7717, 16),
    156 => to_signed(7766, 16),
    157 => to_signed(7815, 16),
    158 => to_signed(7864, 16),
    159 => to_signed(7912, 16),
    160 => to_signed(7961, 16),
    161 => to_signed(8010, 16),
    162 => to_signed(8059, 16),
    163 => to_signed(8107, 16),
    164 => to_signed(8156, 16),
    165 => to_signed(8205, 16),
    166 => to_signed(8253, 16),
    167 => to_signed(8302, 16),
    168 => to_signed(8351, 16),
    169 => to_signed(8399, 16),
    170 => to_signed(8448, 16),
    171 => to_signed(8496, 16),
    172 => to_signed(8545, 16),
    173 => to_signed(8593, 16),
    174 => to_signed(8642, 16),
    175 => to_signed(8690, 16),
    176 => to_signed(8739, 16),
    177 => to_signed(8787, 16),
    178 => to_signed(8836, 16),
    179 => to_signed(8884, 16),
    180 => to_signed(8932, 16),
    181 => to_signed(8981, 16),
    182 => to_signed(9029, 16),
    183 => to_signed(9077, 16),
    184 => to_signed(9126, 16),
    185 => to_signed(9174, 16),
    186 => to_signed(9222, 16),
    187 => to_signed(9270, 16),
    188 => to_signed(9319, 16),
    189 => to_signed(9367, 16),
    190 => to_signed(9415, 16),
    191 => to_signed(9463, 16),
    192 => to_signed(9511, 16),
    193 => to_signed(9559, 16),
    194 => to_signed(9607, 16),
    195 => to_signed(9655, 16),
    196 => to_signed(9703, 16),
    197 => to_signed(9751, 16),
    198 => to_signed(9799, 16),
    199 => to_signed(9847, 16),
    200 => to_signed(9895, 16),
    201 => to_signed(9943, 16),
    202 => to_signed(9991, 16),
    203 => to_signed(10039, 16),
    204 => to_signed(10087, 16),
    205 => to_signed(10135, 16),
    206 => to_signed(10182, 16),
    207 => to_signed(10230, 16),
    208 => to_signed(10278, 16),
    209 => to_signed(10326, 16),
    210 => to_signed(10373, 16),
    211 => to_signed(10421, 16),
    212 => to_signed(10469, 16),
    213 => to_signed(10516, 16),
    214 => to_signed(10564, 16),
    215 => to_signed(10611, 16),
    216 => to_signed(10659, 16),
    217 => to_signed(10706, 16),
    218 => to_signed(10754, 16),
    219 => to_signed(10801, 16),
    220 => to_signed(10849, 16),
    221 => to_signed(10896, 16),
    222 => to_signed(10944, 16),
    223 => to_signed(10991, 16),
    224 => to_signed(11038, 16),
    225 => to_signed(11086, 16),
    226 => to_signed(11133, 16),
    227 => to_signed(11180, 16),
    228 => to_signed(11227, 16),
    229 => to_signed(11275, 16),
    230 => to_signed(11322, 16),
    231 => to_signed(11369, 16),
    232 => to_signed(11416, 16),
    233 => to_signed(11463, 16),
    234 => to_signed(11510, 16),
    235 => to_signed(11557, 16),
    236 => to_signed(11604, 16),
    237 => to_signed(11651, 16),
    238 => to_signed(11698, 16),
    239 => to_signed(11745, 16),
    240 => to_signed(11792, 16),
    241 => to_signed(11839, 16),
    242 => to_signed(11886, 16),
    243 => to_signed(11933, 16),
    244 => to_signed(11980, 16),
    245 => to_signed(12026, 16),
    246 => to_signed(12073, 16),
    247 => to_signed(12120, 16),
    248 => to_signed(12166, 16),
    249 => to_signed(12213, 16),
    250 => to_signed(12260, 16),
    251 => to_signed(12306, 16),
    252 => to_signed(12353, 16),
    253 => to_signed(12399, 16),
    254 => to_signed(12446, 16),
    255 => to_signed(12492, 16),
    256 => to_signed(12539, 16),
    257 => to_signed(12585, 16),
    258 => to_signed(12632, 16),
    259 => to_signed(12678, 16),
    260 => to_signed(12724, 16),
    261 => to_signed(12771, 16),
    262 => to_signed(12817, 16),
    263 => to_signed(12863, 16),
    264 => to_signed(12909, 16),
    265 => to_signed(12956, 16),
    266 => to_signed(13002, 16),
    267 => to_signed(13048, 16),
    268 => to_signed(13094, 16),
    269 => to_signed(13140, 16),
    270 => to_signed(13186, 16),
    271 => to_signed(13232, 16),
    272 => to_signed(13278, 16),
    273 => to_signed(13324, 16),
    274 => to_signed(13370, 16),
    275 => to_signed(13416, 16),
    276 => to_signed(13462, 16),
    277 => to_signed(13507, 16),
    278 => to_signed(13553, 16),
    279 => to_signed(13599, 16),
    280 => to_signed(13645, 16),
    281 => to_signed(13690, 16),
    282 => to_signed(13736, 16),
    283 => to_signed(13782, 16),
    284 => to_signed(13827, 16),
    285 => to_signed(13873, 16),
    286 => to_signed(13918, 16),
    287 => to_signed(13964, 16),
    288 => to_signed(14009, 16),
    289 => to_signed(14055, 16),
    290 => to_signed(14100, 16),
    291 => to_signed(14145, 16),
    292 => to_signed(14191, 16),
    293 => to_signed(14236, 16),
    294 => to_signed(14281, 16),
    295 => to_signed(14326, 16),
    296 => to_signed(14372, 16),
    297 => to_signed(14417, 16),
    298 => to_signed(14462, 16),
    299 => to_signed(14507, 16),
    300 => to_signed(14552, 16),
    301 => to_signed(14597, 16),
    302 => to_signed(14642, 16),
    303 => to_signed(14687, 16),
    304 => to_signed(14732, 16),
    305 => to_signed(14777, 16),
    306 => to_signed(14822, 16),
    307 => to_signed(14866, 16),
    308 => to_signed(14911, 16),
    309 => to_signed(14956, 16),
    310 => to_signed(15001, 16),
    311 => to_signed(15045, 16),
    312 => to_signed(15090, 16),
    313 => to_signed(15135, 16),
    314 => to_signed(15179, 16),
    315 => to_signed(15224, 16),
    316 => to_signed(15268, 16),
    317 => to_signed(15313, 16),
    318 => to_signed(15357, 16),
    319 => to_signed(15401, 16),
    320 => to_signed(15446, 16),
    321 => to_signed(15490, 16),
    322 => to_signed(15534, 16),
    323 => to_signed(15579, 16),
    324 => to_signed(15623, 16),
    325 => to_signed(15667, 16),
    326 => to_signed(15711, 16),
    327 => to_signed(15755, 16),
    328 => to_signed(15799, 16),
    329 => to_signed(15843, 16),
    330 => to_signed(15887, 16),
    331 => to_signed(15931, 16),
    332 => to_signed(15975, 16),
    333 => to_signed(16019, 16),
    334 => to_signed(16063, 16),
    335 => to_signed(16107, 16),
    336 => to_signed(16150, 16),
    337 => to_signed(16194, 16),
    338 => to_signed(16238, 16),
    339 => to_signed(16281, 16),
    340 => to_signed(16325, 16),
    341 => to_signed(16368, 16),
    342 => to_signed(16412, 16),
    343 => to_signed(16455, 16),
    344 => to_signed(16499, 16),
    345 => to_signed(16542, 16),
    346 => to_signed(16586, 16),
    347 => to_signed(16629, 16),
    348 => to_signed(16672, 16),
    349 => to_signed(16716, 16),
    350 => to_signed(16759, 16),
    351 => to_signed(16802, 16),
    352 => to_signed(16845, 16),
    353 => to_signed(16888, 16),
    354 => to_signed(16931, 16),
    355 => to_signed(16974, 16),
    356 => to_signed(17017, 16),
    357 => to_signed(17060, 16),
    358 => to_signed(17103, 16),
    359 => to_signed(17146, 16),
    360 => to_signed(17189, 16),
    361 => to_signed(17232, 16),
    362 => to_signed(17274, 16),
    363 => to_signed(17317, 16),
    364 => to_signed(17360, 16),
    365 => to_signed(17402, 16),
    366 => to_signed(17445, 16),
    367 => to_signed(17487, 16),
    368 => to_signed(17530, 16),
    369 => to_signed(17572, 16),
    370 => to_signed(17615, 16),
    371 => to_signed(17657, 16),
    372 => to_signed(17699, 16),
    373 => to_signed(17742, 16),
    374 => to_signed(17784, 16),
    375 => to_signed(17826, 16),
    376 => to_signed(17868, 16),
    377 => to_signed(17910, 16),
    378 => to_signed(17952, 16),
    379 => to_signed(17994, 16),
    380 => to_signed(18036, 16),
    381 => to_signed(18078, 16),
    382 => to_signed(18120, 16),
    383 => to_signed(18162, 16),
    384 => to_signed(18204, 16),
    385 => to_signed(18246, 16),
    386 => to_signed(18287, 16),
    387 => to_signed(18329, 16),
    388 => to_signed(18371, 16),
    389 => to_signed(18412, 16),
    390 => to_signed(18454, 16),
    391 => to_signed(18495, 16),
    392 => to_signed(18537, 16),
    393 => to_signed(18578, 16),
    394 => to_signed(18620, 16),
    395 => to_signed(18661, 16),
    396 => to_signed(18702, 16),
    397 => to_signed(18744, 16),
    398 => to_signed(18785, 16),
    399 => to_signed(18826, 16),
    400 => to_signed(18867, 16),
    401 => to_signed(18908, 16),
    402 => to_signed(18949, 16),
    403 => to_signed(18990, 16),
    404 => to_signed(19031, 16),
    405 => to_signed(19072, 16),
    406 => to_signed(19113, 16),
    407 => to_signed(19154, 16),
    408 => to_signed(19194, 16),
    409 => to_signed(19235, 16),
    410 => to_signed(19276, 16),
    411 => to_signed(19316, 16),
    412 => to_signed(19357, 16),
    413 => to_signed(19397, 16),
    414 => to_signed(19438, 16),
    415 => to_signed(19478, 16),
    416 => to_signed(19519, 16),
    417 => to_signed(19559, 16),
    418 => to_signed(19599, 16),
    419 => to_signed(19640, 16),
    420 => to_signed(19680, 16),
    421 => to_signed(19720, 16),
    422 => to_signed(19760, 16),
    423 => to_signed(19800, 16),
    424 => to_signed(19840, 16),
    425 => to_signed(19880, 16),
    426 => to_signed(19920, 16),
    427 => to_signed(19960, 16),
    428 => to_signed(20000, 16),
    429 => to_signed(20040, 16),
    430 => to_signed(20079, 16),
    431 => to_signed(20119, 16),
    432 => to_signed(20159, 16),
    433 => to_signed(20198, 16),
    434 => to_signed(20238, 16),
    435 => to_signed(20277, 16),
    436 => to_signed(20317, 16),
    437 => to_signed(20356, 16),
    438 => to_signed(20396, 16),
    439 => to_signed(20435, 16),
    440 => to_signed(20474, 16),
    441 => to_signed(20513, 16),
    442 => to_signed(20553, 16),
    443 => to_signed(20592, 16),
    444 => to_signed(20631, 16),
    445 => to_signed(20670, 16),
    446 => to_signed(20709, 16),
    447 => to_signed(20748, 16),
    448 => to_signed(20787, 16),
    449 => to_signed(20825, 16),
    450 => to_signed(20864, 16),
    451 => to_signed(20903, 16),
    452 => to_signed(20942, 16),
    453 => to_signed(20980, 16),
    454 => to_signed(21019, 16),
    455 => to_signed(21057, 16),
    456 => to_signed(21096, 16),
    457 => to_signed(21134, 16),
    458 => to_signed(21173, 16),
    459 => to_signed(21211, 16),
    460 => to_signed(21249, 16),
    461 => to_signed(21288, 16),
    462 => to_signed(21326, 16),
    463 => to_signed(21364, 16),
    464 => to_signed(21402, 16),
    465 => to_signed(21440, 16),
    466 => to_signed(21478, 16),
    467 => to_signed(21516, 16),
    468 => to_signed(21554, 16),
    469 => to_signed(21592, 16),
    470 => to_signed(21629, 16),
    471 => to_signed(21667, 16),
    472 => to_signed(21705, 16),
    473 => to_signed(21743, 16),
    474 => to_signed(21780, 16),
    475 => to_signed(21818, 16),
    476 => to_signed(21855, 16),
    477 => to_signed(21893, 16),
    478 => to_signed(21930, 16),
    479 => to_signed(21967, 16),
    480 => to_signed(22004, 16),
    481 => to_signed(22042, 16),
    482 => to_signed(22079, 16),
    483 => to_signed(22116, 16),
    484 => to_signed(22153, 16),
    485 => to_signed(22190, 16),
    486 => to_signed(22227, 16),
    487 => to_signed(22264, 16),
    488 => to_signed(22301, 16),
    489 => to_signed(22338, 16),
    490 => to_signed(22374, 16),
    491 => to_signed(22411, 16),
    492 => to_signed(22448, 16),
    493 => to_signed(22484, 16),
    494 => to_signed(22521, 16),
    495 => to_signed(22557, 16),
    496 => to_signed(22594, 16),
    497 => to_signed(22630, 16),
    498 => to_signed(22666, 16),
    499 => to_signed(22703, 16),
    500 => to_signed(22739, 16),
    501 => to_signed(22775, 16),
    502 => to_signed(22811, 16),
    503 => to_signed(22847, 16),
    504 => to_signed(22883, 16),
    505 => to_signed(22919, 16),
    506 => to_signed(22955, 16),
    507 => to_signed(22991, 16),
    508 => to_signed(23027, 16),
    509 => to_signed(23062, 16),
    510 => to_signed(23098, 16),
    511 => to_signed(23134, 16),
    512 => to_signed(23169, 16),
    513 => to_signed(23205, 16),
    514 => to_signed(23240, 16),
    515 => to_signed(23276, 16),
    516 => to_signed(23311, 16),
    517 => to_signed(23346, 16),
    518 => to_signed(23382, 16),
    519 => to_signed(23417, 16),
    520 => to_signed(23452, 16),
    521 => to_signed(23487, 16),
    522 => to_signed(23522, 16),
    523 => to_signed(23557, 16),
    524 => to_signed(23592, 16),
    525 => to_signed(23627, 16),
    526 => to_signed(23661, 16),
    527 => to_signed(23696, 16),
    528 => to_signed(23731, 16),
    529 => to_signed(23766, 16),
    530 => to_signed(23800, 16),
    531 => to_signed(23835, 16),
    532 => to_signed(23869, 16),
    533 => to_signed(23903, 16),
    534 => to_signed(23938, 16),
    535 => to_signed(23972, 16),
    536 => to_signed(24006, 16),
    537 => to_signed(24041, 16),
    538 => to_signed(24075, 16),
    539 => to_signed(24109, 16),
    540 => to_signed(24143, 16),
    541 => to_signed(24177, 16),
    542 => to_signed(24211, 16),
    543 => to_signed(24244, 16),
    544 => to_signed(24278, 16),
    545 => to_signed(24312, 16),
    546 => to_signed(24346, 16),
    547 => to_signed(24379, 16),
    548 => to_signed(24413, 16),
    549 => to_signed(24446, 16),
    550 => to_signed(24480, 16),
    551 => to_signed(24513, 16),
    552 => to_signed(24546, 16),
    553 => to_signed(24580, 16),
    554 => to_signed(24613, 16),
    555 => to_signed(24646, 16),
    556 => to_signed(24679, 16),
    557 => to_signed(24712, 16),
    558 => to_signed(24745, 16),
    559 => to_signed(24778, 16),
    560 => to_signed(24811, 16),
    561 => to_signed(24844, 16),
    562 => to_signed(24877, 16),
    563 => to_signed(24909, 16),
    564 => to_signed(24942, 16),
    565 => to_signed(24974, 16),
    566 => to_signed(25007, 16),
    567 => to_signed(25039, 16),
    568 => to_signed(25072, 16),
    569 => to_signed(25104, 16),
    570 => to_signed(25136, 16),
    571 => to_signed(25169, 16),
    572 => to_signed(25201, 16),
    573 => to_signed(25233, 16),
    574 => to_signed(25265, 16),
    575 => to_signed(25297, 16),
    576 => to_signed(25329, 16),
    577 => to_signed(25361, 16),
    578 => to_signed(25392, 16),
    579 => to_signed(25424, 16),
    580 => to_signed(25456, 16),
    581 => to_signed(25487, 16),
    582 => to_signed(25519, 16),
    583 => to_signed(25550, 16),
    584 => to_signed(25582, 16),
    585 => to_signed(25613, 16),
    586 => to_signed(25645, 16),
    587 => to_signed(25676, 16),
    588 => to_signed(25707, 16),
    589 => to_signed(25738, 16),
    590 => to_signed(25769, 16),
    591 => to_signed(25800, 16),
    592 => to_signed(25831, 16),
    593 => to_signed(25862, 16),
    594 => to_signed(25893, 16),
    595 => to_signed(25924, 16),
    596 => to_signed(25954, 16),
    597 => to_signed(25985, 16),
    598 => to_signed(26016, 16),
    599 => to_signed(26046, 16),
    600 => to_signed(26077, 16),
    601 => to_signed(26107, 16),
    602 => to_signed(26137, 16),
    603 => to_signed(26168, 16),
    604 => to_signed(26198, 16),
    605 => to_signed(26228, 16),
    606 => to_signed(26258, 16),
    607 => to_signed(26288, 16),
    608 => to_signed(26318, 16),
    609 => to_signed(26348, 16),
    610 => to_signed(26378, 16),
    611 => to_signed(26408, 16),
    612 => to_signed(26437, 16),
    613 => to_signed(26467, 16),
    614 => to_signed(26497, 16),
    615 => to_signed(26526, 16),
    616 => to_signed(26556, 16),
    617 => to_signed(26585, 16),
    618 => to_signed(26615, 16),
    619 => to_signed(26644, 16),
    620 => to_signed(26673, 16),
    621 => to_signed(26702, 16),
    622 => to_signed(26731, 16),
    623 => to_signed(26760, 16),
    624 => to_signed(26789, 16),
    625 => to_signed(26818, 16),
    626 => to_signed(26847, 16),
    627 => to_signed(26876, 16),
    628 => to_signed(26905, 16),
    629 => to_signed(26933, 16),
    630 => to_signed(26962, 16),
    631 => to_signed(26990, 16),
    632 => to_signed(27019, 16),
    633 => to_signed(27047, 16),
    634 => to_signed(27076, 16),
    635 => to_signed(27104, 16),
    636 => to_signed(27132, 16),
    637 => to_signed(27160, 16),
    638 => to_signed(27188, 16),
    639 => to_signed(27216, 16),
    640 => to_signed(27244, 16),
    641 => to_signed(27272, 16),
    642 => to_signed(27300, 16),
    643 => to_signed(27328, 16),
    644 => to_signed(27355, 16),
    645 => to_signed(27383, 16),
    646 => to_signed(27411, 16),
    647 => to_signed(27438, 16),
    648 => to_signed(27466, 16),
    649 => to_signed(27493, 16),
    650 => to_signed(27520, 16),
    651 => to_signed(27548, 16),
    652 => to_signed(27575, 16),
    653 => to_signed(27602, 16),
    654 => to_signed(27629, 16),
    655 => to_signed(27656, 16),
    656 => to_signed(27683, 16),
    657 => to_signed(27710, 16),
    658 => to_signed(27736, 16),
    659 => to_signed(27763, 16),
    660 => to_signed(27790, 16),
    661 => to_signed(27816, 16),
    662 => to_signed(27843, 16),
    663 => to_signed(27869, 16),
    664 => to_signed(27896, 16),
    665 => to_signed(27922, 16),
    666 => to_signed(27948, 16),
    667 => to_signed(27975, 16),
    668 => to_signed(28001, 16),
    669 => to_signed(28027, 16),
    670 => to_signed(28053, 16),
    671 => to_signed(28079, 16),
    672 => to_signed(28105, 16),
    673 => to_signed(28131, 16),
    674 => to_signed(28156, 16),
    675 => to_signed(28182, 16),
    676 => to_signed(28208, 16),
    677 => to_signed(28233, 16),
    678 => to_signed(28259, 16),
    679 => to_signed(28284, 16),
    680 => to_signed(28309, 16),
    681 => to_signed(28335, 16),
    682 => to_signed(28360, 16),
    683 => to_signed(28385, 16),
    684 => to_signed(28410, 16),
    685 => to_signed(28435, 16),
    686 => to_signed(28460, 16),
    687 => to_signed(28485, 16),
    688 => to_signed(28510, 16),
    689 => to_signed(28534, 16),
    690 => to_signed(28559, 16),
    691 => to_signed(28584, 16),
    692 => to_signed(28608, 16),
    693 => to_signed(28633, 16),
    694 => to_signed(28657, 16),
    695 => to_signed(28681, 16),
    696 => to_signed(28706, 16),
    697 => to_signed(28730, 16),
    698 => to_signed(28754, 16),
    699 => to_signed(28778, 16),
    700 => to_signed(28802, 16),
    701 => to_signed(28826, 16),
    702 => to_signed(28850, 16),
    703 => to_signed(28874, 16),
    704 => to_signed(28897, 16),
    705 => to_signed(28921, 16),
    706 => to_signed(28945, 16),
    707 => to_signed(28968, 16),
    708 => to_signed(28992, 16),
    709 => to_signed(29015, 16),
    710 => to_signed(29038, 16),
    711 => to_signed(29062, 16),
    712 => to_signed(29085, 16),
    713 => to_signed(29108, 16),
    714 => to_signed(29131, 16),
    715 => to_signed(29154, 16),
    716 => to_signed(29177, 16),
    717 => to_signed(29200, 16),
    718 => to_signed(29222, 16),
    719 => to_signed(29245, 16),
    720 => to_signed(29268, 16),
    721 => to_signed(29290, 16),
    722 => to_signed(29313, 16),
    723 => to_signed(29335, 16),
    724 => to_signed(29358, 16),
    725 => to_signed(29380, 16),
    726 => to_signed(29402, 16),
    727 => to_signed(29424, 16),
    728 => to_signed(29446, 16),
    729 => to_signed(29468, 16),
    730 => to_signed(29490, 16),
    731 => to_signed(29512, 16),
    732 => to_signed(29534, 16),
    733 => to_signed(29556, 16),
    734 => to_signed(29577, 16),
    735 => to_signed(29599, 16),
    736 => to_signed(29621, 16),
    737 => to_signed(29642, 16),
    738 => to_signed(29663, 16),
    739 => to_signed(29685, 16),
    740 => to_signed(29706, 16),
    741 => to_signed(29727, 16),
    742 => to_signed(29748, 16),
    743 => to_signed(29769, 16),
    744 => to_signed(29790, 16),
    745 => to_signed(29811, 16),
    746 => to_signed(29832, 16),
    747 => to_signed(29853, 16),
    748 => to_signed(29873, 16),
    749 => to_signed(29894, 16),
    750 => to_signed(29915, 16),
    751 => to_signed(29935, 16),
    752 => to_signed(29955, 16),
    753 => to_signed(29976, 16),
    754 => to_signed(29996, 16),
    755 => to_signed(30016, 16),
    756 => to_signed(30036, 16),
    757 => to_signed(30056, 16),
    758 => to_signed(30076, 16),
    759 => to_signed(30096, 16),
    760 => to_signed(30116, 16),
    761 => to_signed(30136, 16),
    762 => to_signed(30156, 16),
    763 => to_signed(30175, 16),
    764 => to_signed(30195, 16),
    765 => to_signed(30214, 16),
    766 => to_signed(30234, 16),
    767 => to_signed(30253, 16),
    768 => to_signed(30272, 16),
    769 => to_signed(30291, 16),
    770 => to_signed(30311, 16),
    771 => to_signed(30330, 16),
    772 => to_signed(30349, 16),
    773 => to_signed(30368, 16),
    774 => to_signed(30386, 16),
    775 => to_signed(30405, 16),
    776 => to_signed(30424, 16),
    777 => to_signed(30442, 16),
    778 => to_signed(30461, 16),
    779 => to_signed(30480, 16),
    780 => to_signed(30498, 16),
    781 => to_signed(30516, 16),
    782 => to_signed(30535, 16),
    783 => to_signed(30553, 16),
    784 => to_signed(30571, 16),
    785 => to_signed(30589, 16),
    786 => to_signed(30607, 16),
    787 => to_signed(30625, 16),
    788 => to_signed(30643, 16),
    789 => to_signed(30660, 16),
    790 => to_signed(30678, 16),
    791 => to_signed(30696, 16),
    792 => to_signed(30713, 16),
    793 => to_signed(30731, 16),
    794 => to_signed(30748, 16),
    795 => to_signed(30766, 16),
    796 => to_signed(30783, 16),
    797 => to_signed(30800, 16),
    798 => to_signed(30817, 16),
    799 => to_signed(30834, 16),
    800 => to_signed(30851, 16),
    801 => to_signed(30868, 16),
    802 => to_signed(30885, 16),
    803 => to_signed(30902, 16),
    804 => to_signed(30918, 16),
    805 => to_signed(30935, 16),
    806 => to_signed(30951, 16),
    807 => to_signed(30968, 16),
    808 => to_signed(30984, 16),
    809 => to_signed(31001, 16),
    810 => to_signed(31017, 16),
    811 => to_signed(31033, 16),
    812 => to_signed(31049, 16),
    813 => to_signed(31065, 16),
    814 => to_signed(31081, 16),
    815 => to_signed(31097, 16),
    816 => to_signed(31113, 16),
    817 => to_signed(31128, 16),
    818 => to_signed(31144, 16),
    819 => to_signed(31160, 16),
    820 => to_signed(31175, 16),
    821 => to_signed(31191, 16),
    822 => to_signed(31206, 16),
    823 => to_signed(31221, 16),
    824 => to_signed(31236, 16),
    825 => to_signed(31252, 16),
    826 => to_signed(31267, 16),
    827 => to_signed(31282, 16),
    828 => to_signed(31297, 16),
    829 => to_signed(31311, 16),
    830 => to_signed(31326, 16),
    831 => to_signed(31341, 16),
    832 => to_signed(31356, 16),
    833 => to_signed(31370, 16),
    834 => to_signed(31385, 16),
    835 => to_signed(31399, 16),
    836 => to_signed(31413, 16),
    837 => to_signed(31428, 16),
    838 => to_signed(31442, 16),
    839 => to_signed(31456, 16),
    840 => to_signed(31470, 16),
    841 => to_signed(31484, 16),
    842 => to_signed(31498, 16),
    843 => to_signed(31512, 16),
    844 => to_signed(31525, 16),
    845 => to_signed(31539, 16),
    846 => to_signed(31553, 16),
    847 => to_signed(31566, 16),
    848 => to_signed(31580, 16),
    849 => to_signed(31593, 16),
    850 => to_signed(31606, 16),
    851 => to_signed(31619, 16),
    852 => to_signed(31633, 16),
    853 => to_signed(31646, 16),
    854 => to_signed(31659, 16),
    855 => to_signed(31672, 16),
    856 => to_signed(31684, 16),
    857 => to_signed(31697, 16),
    858 => to_signed(31710, 16),
    859 => to_signed(31723, 16),
    860 => to_signed(31735, 16),
    861 => to_signed(31748, 16),
    862 => to_signed(31760, 16),
    863 => to_signed(31772, 16),
    864 => to_signed(31785, 16),
    865 => to_signed(31797, 16),
    866 => to_signed(31809, 16),
    867 => to_signed(31821, 16),
    868 => to_signed(31833, 16),
    869 => to_signed(31845, 16),
    870 => to_signed(31856, 16),
    871 => to_signed(31868, 16),
    872 => to_signed(31880, 16),
    873 => to_signed(31891, 16),
    874 => to_signed(31903, 16),
    875 => to_signed(31914, 16),
    876 => to_signed(31926, 16),
    877 => to_signed(31937, 16),
    878 => to_signed(31948, 16),
    879 => to_signed(31959, 16),
    880 => to_signed(31970, 16),
    881 => to_signed(31981, 16),
    882 => to_signed(31992, 16),
    883 => to_signed(32003, 16),
    884 => to_signed(32014, 16),
    885 => to_signed(32024, 16),
    886 => to_signed(32035, 16),
    887 => to_signed(32046, 16),
    888 => to_signed(32056, 16),
    889 => to_signed(32066, 16),
    890 => to_signed(32077, 16),
    891 => to_signed(32087, 16),
    892 => to_signed(32097, 16),
    893 => to_signed(32107, 16),
    894 => to_signed(32117, 16),
    895 => to_signed(32127, 16),
    896 => to_signed(32137, 16),
    897 => to_signed(32147, 16),
    898 => to_signed(32156, 16),
    899 => to_signed(32166, 16),
    900 => to_signed(32176, 16),
    901 => to_signed(32185, 16),
    902 => to_signed(32194, 16),
    903 => to_signed(32204, 16),
    904 => to_signed(32213, 16),
    905 => to_signed(32222, 16),
    906 => to_signed(32231, 16),
    907 => to_signed(32240, 16),
    908 => to_signed(32249, 16),
    909 => to_signed(32258, 16),
    910 => to_signed(32267, 16),
    911 => to_signed(32275, 16),
    912 => to_signed(32284, 16),
    913 => to_signed(32293, 16),
    914 => to_signed(32301, 16),
    915 => to_signed(32310, 16),
    916 => to_signed(32318, 16),
    917 => to_signed(32326, 16),
    918 => to_signed(32334, 16),
    919 => to_signed(32342, 16),
    920 => to_signed(32350, 16),
    921 => to_signed(32358, 16),
    922 => to_signed(32366, 16),
    923 => to_signed(32374, 16),
    924 => to_signed(32382, 16),
    925 => to_signed(32389, 16),
    926 => to_signed(32397, 16),
    927 => to_signed(32404, 16),
    928 => to_signed(32412, 16),
    929 => to_signed(32419, 16),
    930 => to_signed(32426, 16),
    931 => to_signed(32434, 16),
    932 => to_signed(32441, 16),
    933 => to_signed(32448, 16),
    934 => to_signed(32455, 16),
    935 => to_signed(32462, 16),
    936 => to_signed(32468, 16),
    937 => to_signed(32475, 16),
    938 => to_signed(32482, 16),
    939 => to_signed(32488, 16),
    940 => to_signed(32495, 16),
    941 => to_signed(32501, 16),
    942 => to_signed(32508, 16),
    943 => to_signed(32514, 16),
    944 => to_signed(32520, 16),
    945 => to_signed(32526, 16),
    946 => to_signed(32532, 16),
    947 => to_signed(32538, 16),
    948 => to_signed(32544, 16),
    949 => to_signed(32550, 16),
    950 => to_signed(32556, 16),
    951 => to_signed(32561, 16),
    952 => to_signed(32567, 16),
    953 => to_signed(32572, 16),
    954 => to_signed(32578, 16),
    955 => to_signed(32583, 16),
    956 => to_signed(32588, 16),
    957 => to_signed(32594, 16),
    958 => to_signed(32599, 16),
    959 => to_signed(32604, 16),
    960 => to_signed(32609, 16),
    961 => to_signed(32614, 16),
    962 => to_signed(32618, 16),
    963 => to_signed(32623, 16),
    964 => to_signed(32628, 16),
    965 => to_signed(32632, 16),
    966 => to_signed(32637, 16),
    967 => to_signed(32641, 16),
    968 => to_signed(32646, 16),
    969 => to_signed(32650, 16),
    970 => to_signed(32654, 16),
    971 => to_signed(32658, 16),
    972 => to_signed(32662, 16),
    973 => to_signed(32666, 16),
    974 => to_signed(32670, 16),
    975 => to_signed(32674, 16),
    976 => to_signed(32678, 16),
    977 => to_signed(32681, 16),
    978 => to_signed(32685, 16),
    979 => to_signed(32688, 16),
    980 => to_signed(32692, 16),
    981 => to_signed(32695, 16),
    982 => to_signed(32699, 16),
    983 => to_signed(32702, 16),
    984 => to_signed(32705, 16),
    985 => to_signed(32708, 16),
    986 => to_signed(32711, 16),
    987 => to_signed(32714, 16),
    988 => to_signed(32717, 16),
    989 => to_signed(32719, 16),
    990 => to_signed(32722, 16),
    991 => to_signed(32725, 16),
    992 => to_signed(32727, 16),
    993 => to_signed(32729, 16),
    994 => to_signed(32732, 16),
    995 => to_signed(32734, 16),
    996 => to_signed(32736, 16),
    997 => to_signed(32738, 16),
    998 => to_signed(32740, 16),
    999 => to_signed(32742, 16),
    1000 => to_signed(32744, 16),
    1001 => to_signed(32746, 16),
    1002 => to_signed(32748, 16),
    1003 => to_signed(32750, 16),
    1004 => to_signed(32751, 16),
    1005 => to_signed(32753, 16),
    1006 => to_signed(32754, 16),
    1007 => to_signed(32755, 16),
    1008 => to_signed(32757, 16),
    1009 => to_signed(32758, 16),
    1010 => to_signed(32759, 16),
    1011 => to_signed(32760, 16),
    1012 => to_signed(32761, 16),
    1013 => to_signed(32762, 16),
    1014 => to_signed(32763, 16),
    1015 => to_signed(32763, 16),
    1016 => to_signed(32764, 16),
    1017 => to_signed(32765, 16),
    1018 => to_signed(32765, 16),
    1019 => to_signed(32766, 16),
    1020 => to_signed(32766, 16),
    1021 => to_signed(32766, 16),
    1022 => to_signed(32766, 16),
    1023 => to_signed(32766, 16),
    1024 => to_signed(32767, 16),
    1025 => to_signed(32766, 16),
    1026 => to_signed(32766, 16),
    1027 => to_signed(32766, 16),
    1028 => to_signed(32766, 16),
    1029 => to_signed(32766, 16),
    1030 => to_signed(32765, 16),
    1031 => to_signed(32765, 16),
    1032 => to_signed(32764, 16),
    1033 => to_signed(32763, 16),
    1034 => to_signed(32763, 16),
    1035 => to_signed(32762, 16),
    1036 => to_signed(32761, 16),
    1037 => to_signed(32760, 16),
    1038 => to_signed(32759, 16),
    1039 => to_signed(32758, 16),
    1040 => to_signed(32757, 16),
    1041 => to_signed(32755, 16),
    1042 => to_signed(32754, 16),
    1043 => to_signed(32753, 16),
    1044 => to_signed(32751, 16),
    1045 => to_signed(32750, 16),
    1046 => to_signed(32748, 16),
    1047 => to_signed(32746, 16),
    1048 => to_signed(32744, 16),
    1049 => to_signed(32742, 16),
    1050 => to_signed(32740, 16),
    1051 => to_signed(32738, 16),
    1052 => to_signed(32736, 16),
    1053 => to_signed(32734, 16),
    1054 => to_signed(32732, 16),
    1055 => to_signed(32729, 16),
    1056 => to_signed(32727, 16),
    1057 => to_signed(32725, 16),
    1058 => to_signed(32722, 16),
    1059 => to_signed(32719, 16),
    1060 => to_signed(32717, 16),
    1061 => to_signed(32714, 16),
    1062 => to_signed(32711, 16),
    1063 => to_signed(32708, 16),
    1064 => to_signed(32705, 16),
    1065 => to_signed(32702, 16),
    1066 => to_signed(32699, 16),
    1067 => to_signed(32695, 16),
    1068 => to_signed(32692, 16),
    1069 => to_signed(32688, 16),
    1070 => to_signed(32685, 16),
    1071 => to_signed(32681, 16),
    1072 => to_signed(32678, 16),
    1073 => to_signed(32674, 16),
    1074 => to_signed(32670, 16),
    1075 => to_signed(32666, 16),
    1076 => to_signed(32662, 16),
    1077 => to_signed(32658, 16),
    1078 => to_signed(32654, 16),
    1079 => to_signed(32650, 16),
    1080 => to_signed(32646, 16),
    1081 => to_signed(32641, 16),
    1082 => to_signed(32637, 16),
    1083 => to_signed(32632, 16),
    1084 => to_signed(32628, 16),
    1085 => to_signed(32623, 16),
    1086 => to_signed(32618, 16),
    1087 => to_signed(32614, 16),
    1088 => to_signed(32609, 16),
    1089 => to_signed(32604, 16),
    1090 => to_signed(32599, 16),
    1091 => to_signed(32594, 16),
    1092 => to_signed(32588, 16),
    1093 => to_signed(32583, 16),
    1094 => to_signed(32578, 16),
    1095 => to_signed(32572, 16),
    1096 => to_signed(32567, 16),
    1097 => to_signed(32561, 16),
    1098 => to_signed(32556, 16),
    1099 => to_signed(32550, 16),
    1100 => to_signed(32544, 16),
    1101 => to_signed(32538, 16),
    1102 => to_signed(32532, 16),
    1103 => to_signed(32526, 16),
    1104 => to_signed(32520, 16),
    1105 => to_signed(32514, 16),
    1106 => to_signed(32508, 16),
    1107 => to_signed(32501, 16),
    1108 => to_signed(32495, 16),
    1109 => to_signed(32488, 16),
    1110 => to_signed(32482, 16),
    1111 => to_signed(32475, 16),
    1112 => to_signed(32468, 16),
    1113 => to_signed(32462, 16),
    1114 => to_signed(32455, 16),
    1115 => to_signed(32448, 16),
    1116 => to_signed(32441, 16),
    1117 => to_signed(32434, 16),
    1118 => to_signed(32426, 16),
    1119 => to_signed(32419, 16),
    1120 => to_signed(32412, 16),
    1121 => to_signed(32404, 16),
    1122 => to_signed(32397, 16),
    1123 => to_signed(32389, 16),
    1124 => to_signed(32382, 16),
    1125 => to_signed(32374, 16),
    1126 => to_signed(32366, 16),
    1127 => to_signed(32358, 16),
    1128 => to_signed(32350, 16),
    1129 => to_signed(32342, 16),
    1130 => to_signed(32334, 16),
    1131 => to_signed(32326, 16),
    1132 => to_signed(32318, 16),
    1133 => to_signed(32310, 16),
    1134 => to_signed(32301, 16),
    1135 => to_signed(32293, 16),
    1136 => to_signed(32284, 16),
    1137 => to_signed(32275, 16),
    1138 => to_signed(32267, 16),
    1139 => to_signed(32258, 16),
    1140 => to_signed(32249, 16),
    1141 => to_signed(32240, 16),
    1142 => to_signed(32231, 16),
    1143 => to_signed(32222, 16),
    1144 => to_signed(32213, 16),
    1145 => to_signed(32204, 16),
    1146 => to_signed(32194, 16),
    1147 => to_signed(32185, 16),
    1148 => to_signed(32176, 16),
    1149 => to_signed(32166, 16),
    1150 => to_signed(32156, 16),
    1151 => to_signed(32147, 16),
    1152 => to_signed(32137, 16),
    1153 => to_signed(32127, 16),
    1154 => to_signed(32117, 16),
    1155 => to_signed(32107, 16),
    1156 => to_signed(32097, 16),
    1157 => to_signed(32087, 16),
    1158 => to_signed(32077, 16),
    1159 => to_signed(32066, 16),
    1160 => to_signed(32056, 16),
    1161 => to_signed(32046, 16),
    1162 => to_signed(32035, 16),
    1163 => to_signed(32024, 16),
    1164 => to_signed(32014, 16),
    1165 => to_signed(32003, 16),
    1166 => to_signed(31992, 16),
    1167 => to_signed(31981, 16),
    1168 => to_signed(31970, 16),
    1169 => to_signed(31959, 16),
    1170 => to_signed(31948, 16),
    1171 => to_signed(31937, 16),
    1172 => to_signed(31926, 16),
    1173 => to_signed(31914, 16),
    1174 => to_signed(31903, 16),
    1175 => to_signed(31891, 16),
    1176 => to_signed(31880, 16),
    1177 => to_signed(31868, 16),
    1178 => to_signed(31856, 16),
    1179 => to_signed(31845, 16),
    1180 => to_signed(31833, 16),
    1181 => to_signed(31821, 16),
    1182 => to_signed(31809, 16),
    1183 => to_signed(31797, 16),
    1184 => to_signed(31785, 16),
    1185 => to_signed(31772, 16),
    1186 => to_signed(31760, 16),
    1187 => to_signed(31748, 16),
    1188 => to_signed(31735, 16),
    1189 => to_signed(31723, 16),
    1190 => to_signed(31710, 16),
    1191 => to_signed(31697, 16),
    1192 => to_signed(31684, 16),
    1193 => to_signed(31672, 16),
    1194 => to_signed(31659, 16),
    1195 => to_signed(31646, 16),
    1196 => to_signed(31633, 16),
    1197 => to_signed(31619, 16),
    1198 => to_signed(31606, 16),
    1199 => to_signed(31593, 16),
    1200 => to_signed(31580, 16),
    1201 => to_signed(31566, 16),
    1202 => to_signed(31553, 16),
    1203 => to_signed(31539, 16),
    1204 => to_signed(31525, 16),
    1205 => to_signed(31512, 16),
    1206 => to_signed(31498, 16),
    1207 => to_signed(31484, 16),
    1208 => to_signed(31470, 16),
    1209 => to_signed(31456, 16),
    1210 => to_signed(31442, 16),
    1211 => to_signed(31428, 16),
    1212 => to_signed(31413, 16),
    1213 => to_signed(31399, 16),
    1214 => to_signed(31385, 16),
    1215 => to_signed(31370, 16),
    1216 => to_signed(31356, 16),
    1217 => to_signed(31341, 16),
    1218 => to_signed(31326, 16),
    1219 => to_signed(31311, 16),
    1220 => to_signed(31297, 16),
    1221 => to_signed(31282, 16),
    1222 => to_signed(31267, 16),
    1223 => to_signed(31252, 16),
    1224 => to_signed(31236, 16),
    1225 => to_signed(31221, 16),
    1226 => to_signed(31206, 16),
    1227 => to_signed(31191, 16),
    1228 => to_signed(31175, 16),
    1229 => to_signed(31160, 16),
    1230 => to_signed(31144, 16),
    1231 => to_signed(31128, 16),
    1232 => to_signed(31113, 16),
    1233 => to_signed(31097, 16),
    1234 => to_signed(31081, 16),
    1235 => to_signed(31065, 16),
    1236 => to_signed(31049, 16),
    1237 => to_signed(31033, 16),
    1238 => to_signed(31017, 16),
    1239 => to_signed(31001, 16),
    1240 => to_signed(30984, 16),
    1241 => to_signed(30968, 16),
    1242 => to_signed(30951, 16),
    1243 => to_signed(30935, 16),
    1244 => to_signed(30918, 16),
    1245 => to_signed(30902, 16),
    1246 => to_signed(30885, 16),
    1247 => to_signed(30868, 16),
    1248 => to_signed(30851, 16),
    1249 => to_signed(30834, 16),
    1250 => to_signed(30817, 16),
    1251 => to_signed(30800, 16),
    1252 => to_signed(30783, 16),
    1253 => to_signed(30766, 16),
    1254 => to_signed(30748, 16),
    1255 => to_signed(30731, 16),
    1256 => to_signed(30713, 16),
    1257 => to_signed(30696, 16),
    1258 => to_signed(30678, 16),
    1259 => to_signed(30660, 16),
    1260 => to_signed(30643, 16),
    1261 => to_signed(30625, 16),
    1262 => to_signed(30607, 16),
    1263 => to_signed(30589, 16),
    1264 => to_signed(30571, 16),
    1265 => to_signed(30553, 16),
    1266 => to_signed(30535, 16),
    1267 => to_signed(30516, 16),
    1268 => to_signed(30498, 16),
    1269 => to_signed(30480, 16),
    1270 => to_signed(30461, 16),
    1271 => to_signed(30442, 16),
    1272 => to_signed(30424, 16),
    1273 => to_signed(30405, 16),
    1274 => to_signed(30386, 16),
    1275 => to_signed(30368, 16),
    1276 => to_signed(30349, 16),
    1277 => to_signed(30330, 16),
    1278 => to_signed(30311, 16),
    1279 => to_signed(30291, 16),
    1280 => to_signed(30272, 16),
    1281 => to_signed(30253, 16),
    1282 => to_signed(30234, 16),
    1283 => to_signed(30214, 16),
    1284 => to_signed(30195, 16),
    1285 => to_signed(30175, 16),
    1286 => to_signed(30156, 16),
    1287 => to_signed(30136, 16),
    1288 => to_signed(30116, 16),
    1289 => to_signed(30096, 16),
    1290 => to_signed(30076, 16),
    1291 => to_signed(30056, 16),
    1292 => to_signed(30036, 16),
    1293 => to_signed(30016, 16),
    1294 => to_signed(29996, 16),
    1295 => to_signed(29976, 16),
    1296 => to_signed(29955, 16),
    1297 => to_signed(29935, 16),
    1298 => to_signed(29915, 16),
    1299 => to_signed(29894, 16),
    1300 => to_signed(29873, 16),
    1301 => to_signed(29853, 16),
    1302 => to_signed(29832, 16),
    1303 => to_signed(29811, 16),
    1304 => to_signed(29790, 16),
    1305 => to_signed(29769, 16),
    1306 => to_signed(29748, 16),
    1307 => to_signed(29727, 16),
    1308 => to_signed(29706, 16),
    1309 => to_signed(29685, 16),
    1310 => to_signed(29663, 16),
    1311 => to_signed(29642, 16),
    1312 => to_signed(29621, 16),
    1313 => to_signed(29599, 16),
    1314 => to_signed(29577, 16),
    1315 => to_signed(29556, 16),
    1316 => to_signed(29534, 16),
    1317 => to_signed(29512, 16),
    1318 => to_signed(29490, 16),
    1319 => to_signed(29468, 16),
    1320 => to_signed(29446, 16),
    1321 => to_signed(29424, 16),
    1322 => to_signed(29402, 16),
    1323 => to_signed(29380, 16),
    1324 => to_signed(29358, 16),
    1325 => to_signed(29335, 16),
    1326 => to_signed(29313, 16),
    1327 => to_signed(29290, 16),
    1328 => to_signed(29268, 16),
    1329 => to_signed(29245, 16),
    1330 => to_signed(29222, 16),
    1331 => to_signed(29200, 16),
    1332 => to_signed(29177, 16),
    1333 => to_signed(29154, 16),
    1334 => to_signed(29131, 16),
    1335 => to_signed(29108, 16),
    1336 => to_signed(29085, 16),
    1337 => to_signed(29062, 16),
    1338 => to_signed(29038, 16),
    1339 => to_signed(29015, 16),
    1340 => to_signed(28992, 16),
    1341 => to_signed(28968, 16),
    1342 => to_signed(28945, 16),
    1343 => to_signed(28921, 16),
    1344 => to_signed(28897, 16),
    1345 => to_signed(28874, 16),
    1346 => to_signed(28850, 16),
    1347 => to_signed(28826, 16),
    1348 => to_signed(28802, 16),
    1349 => to_signed(28778, 16),
    1350 => to_signed(28754, 16),
    1351 => to_signed(28730, 16),
    1352 => to_signed(28706, 16),
    1353 => to_signed(28681, 16),
    1354 => to_signed(28657, 16),
    1355 => to_signed(28633, 16),
    1356 => to_signed(28608, 16),
    1357 => to_signed(28584, 16),
    1358 => to_signed(28559, 16),
    1359 => to_signed(28534, 16),
    1360 => to_signed(28510, 16),
    1361 => to_signed(28485, 16),
    1362 => to_signed(28460, 16),
    1363 => to_signed(28435, 16),
    1364 => to_signed(28410, 16),
    1365 => to_signed(28385, 16),
    1366 => to_signed(28360, 16),
    1367 => to_signed(28335, 16),
    1368 => to_signed(28309, 16),
    1369 => to_signed(28284, 16),
    1370 => to_signed(28259, 16),
    1371 => to_signed(28233, 16),
    1372 => to_signed(28208, 16),
    1373 => to_signed(28182, 16),
    1374 => to_signed(28156, 16),
    1375 => to_signed(28131, 16),
    1376 => to_signed(28105, 16),
    1377 => to_signed(28079, 16),
    1378 => to_signed(28053, 16),
    1379 => to_signed(28027, 16),
    1380 => to_signed(28001, 16),
    1381 => to_signed(27975, 16),
    1382 => to_signed(27948, 16),
    1383 => to_signed(27922, 16),
    1384 => to_signed(27896, 16),
    1385 => to_signed(27869, 16),
    1386 => to_signed(27843, 16),
    1387 => to_signed(27816, 16),
    1388 => to_signed(27790, 16),
    1389 => to_signed(27763, 16),
    1390 => to_signed(27736, 16),
    1391 => to_signed(27710, 16),
    1392 => to_signed(27683, 16),
    1393 => to_signed(27656, 16),
    1394 => to_signed(27629, 16),
    1395 => to_signed(27602, 16),
    1396 => to_signed(27575, 16),
    1397 => to_signed(27548, 16),
    1398 => to_signed(27520, 16),
    1399 => to_signed(27493, 16),
    1400 => to_signed(27466, 16),
    1401 => to_signed(27438, 16),
    1402 => to_signed(27411, 16),
    1403 => to_signed(27383, 16),
    1404 => to_signed(27355, 16),
    1405 => to_signed(27328, 16),
    1406 => to_signed(27300, 16),
    1407 => to_signed(27272, 16),
    1408 => to_signed(27244, 16),
    1409 => to_signed(27216, 16),
    1410 => to_signed(27188, 16),
    1411 => to_signed(27160, 16),
    1412 => to_signed(27132, 16),
    1413 => to_signed(27104, 16),
    1414 => to_signed(27076, 16),
    1415 => to_signed(27047, 16),
    1416 => to_signed(27019, 16),
    1417 => to_signed(26990, 16),
    1418 => to_signed(26962, 16),
    1419 => to_signed(26933, 16),
    1420 => to_signed(26905, 16),
    1421 => to_signed(26876, 16),
    1422 => to_signed(26847, 16),
    1423 => to_signed(26818, 16),
    1424 => to_signed(26789, 16),
    1425 => to_signed(26760, 16),
    1426 => to_signed(26731, 16),
    1427 => to_signed(26702, 16),
    1428 => to_signed(26673, 16),
    1429 => to_signed(26644, 16),
    1430 => to_signed(26615, 16),
    1431 => to_signed(26585, 16),
    1432 => to_signed(26556, 16),
    1433 => to_signed(26526, 16),
    1434 => to_signed(26497, 16),
    1435 => to_signed(26467, 16),
    1436 => to_signed(26437, 16),
    1437 => to_signed(26408, 16),
    1438 => to_signed(26378, 16),
    1439 => to_signed(26348, 16),
    1440 => to_signed(26318, 16),
    1441 => to_signed(26288, 16),
    1442 => to_signed(26258, 16),
    1443 => to_signed(26228, 16),
    1444 => to_signed(26198, 16),
    1445 => to_signed(26168, 16),
    1446 => to_signed(26137, 16),
    1447 => to_signed(26107, 16),
    1448 => to_signed(26077, 16),
    1449 => to_signed(26046, 16),
    1450 => to_signed(26016, 16),
    1451 => to_signed(25985, 16),
    1452 => to_signed(25954, 16),
    1453 => to_signed(25924, 16),
    1454 => to_signed(25893, 16),
    1455 => to_signed(25862, 16),
    1456 => to_signed(25831, 16),
    1457 => to_signed(25800, 16),
    1458 => to_signed(25769, 16),
    1459 => to_signed(25738, 16),
    1460 => to_signed(25707, 16),
    1461 => to_signed(25676, 16),
    1462 => to_signed(25645, 16),
    1463 => to_signed(25613, 16),
    1464 => to_signed(25582, 16),
    1465 => to_signed(25550, 16),
    1466 => to_signed(25519, 16),
    1467 => to_signed(25487, 16),
    1468 => to_signed(25456, 16),
    1469 => to_signed(25424, 16),
    1470 => to_signed(25392, 16),
    1471 => to_signed(25361, 16),
    1472 => to_signed(25329, 16),
    1473 => to_signed(25297, 16),
    1474 => to_signed(25265, 16),
    1475 => to_signed(25233, 16),
    1476 => to_signed(25201, 16),
    1477 => to_signed(25169, 16),
    1478 => to_signed(25136, 16),
    1479 => to_signed(25104, 16),
    1480 => to_signed(25072, 16),
    1481 => to_signed(25039, 16),
    1482 => to_signed(25007, 16),
    1483 => to_signed(24974, 16),
    1484 => to_signed(24942, 16),
    1485 => to_signed(24909, 16),
    1486 => to_signed(24877, 16),
    1487 => to_signed(24844, 16),
    1488 => to_signed(24811, 16),
    1489 => to_signed(24778, 16),
    1490 => to_signed(24745, 16),
    1491 => to_signed(24712, 16),
    1492 => to_signed(24679, 16),
    1493 => to_signed(24646, 16),
    1494 => to_signed(24613, 16),
    1495 => to_signed(24580, 16),
    1496 => to_signed(24546, 16),
    1497 => to_signed(24513, 16),
    1498 => to_signed(24480, 16),
    1499 => to_signed(24446, 16),
    1500 => to_signed(24413, 16),
    1501 => to_signed(24379, 16),
    1502 => to_signed(24346, 16),
    1503 => to_signed(24312, 16),
    1504 => to_signed(24278, 16),
    1505 => to_signed(24244, 16),
    1506 => to_signed(24211, 16),
    1507 => to_signed(24177, 16),
    1508 => to_signed(24143, 16),
    1509 => to_signed(24109, 16),
    1510 => to_signed(24075, 16),
    1511 => to_signed(24041, 16),
    1512 => to_signed(24006, 16),
    1513 => to_signed(23972, 16),
    1514 => to_signed(23938, 16),
    1515 => to_signed(23903, 16),
    1516 => to_signed(23869, 16),
    1517 => to_signed(23835, 16),
    1518 => to_signed(23800, 16),
    1519 => to_signed(23766, 16),
    1520 => to_signed(23731, 16),
    1521 => to_signed(23696, 16),
    1522 => to_signed(23661, 16),
    1523 => to_signed(23627, 16),
    1524 => to_signed(23592, 16),
    1525 => to_signed(23557, 16),
    1526 => to_signed(23522, 16),
    1527 => to_signed(23487, 16),
    1528 => to_signed(23452, 16),
    1529 => to_signed(23417, 16),
    1530 => to_signed(23382, 16),
    1531 => to_signed(23346, 16),
    1532 => to_signed(23311, 16),
    1533 => to_signed(23276, 16),
    1534 => to_signed(23240, 16),
    1535 => to_signed(23205, 16),
    1536 => to_signed(23169, 16),
    1537 => to_signed(23134, 16),
    1538 => to_signed(23098, 16),
    1539 => to_signed(23062, 16),
    1540 => to_signed(23027, 16),
    1541 => to_signed(22991, 16),
    1542 => to_signed(22955, 16),
    1543 => to_signed(22919, 16),
    1544 => to_signed(22883, 16),
    1545 => to_signed(22847, 16),
    1546 => to_signed(22811, 16),
    1547 => to_signed(22775, 16),
    1548 => to_signed(22739, 16),
    1549 => to_signed(22703, 16),
    1550 => to_signed(22666, 16),
    1551 => to_signed(22630, 16),
    1552 => to_signed(22594, 16),
    1553 => to_signed(22557, 16),
    1554 => to_signed(22521, 16),
    1555 => to_signed(22484, 16),
    1556 => to_signed(22448, 16),
    1557 => to_signed(22411, 16),
    1558 => to_signed(22374, 16),
    1559 => to_signed(22338, 16),
    1560 => to_signed(22301, 16),
    1561 => to_signed(22264, 16),
    1562 => to_signed(22227, 16),
    1563 => to_signed(22190, 16),
    1564 => to_signed(22153, 16),
    1565 => to_signed(22116, 16),
    1566 => to_signed(22079, 16),
    1567 => to_signed(22042, 16),
    1568 => to_signed(22004, 16),
    1569 => to_signed(21967, 16),
    1570 => to_signed(21930, 16),
    1571 => to_signed(21893, 16),
    1572 => to_signed(21855, 16),
    1573 => to_signed(21818, 16),
    1574 => to_signed(21780, 16),
    1575 => to_signed(21743, 16),
    1576 => to_signed(21705, 16),
    1577 => to_signed(21667, 16),
    1578 => to_signed(21629, 16),
    1579 => to_signed(21592, 16),
    1580 => to_signed(21554, 16),
    1581 => to_signed(21516, 16),
    1582 => to_signed(21478, 16),
    1583 => to_signed(21440, 16),
    1584 => to_signed(21402, 16),
    1585 => to_signed(21364, 16),
    1586 => to_signed(21326, 16),
    1587 => to_signed(21288, 16),
    1588 => to_signed(21249, 16),
    1589 => to_signed(21211, 16),
    1590 => to_signed(21173, 16),
    1591 => to_signed(21134, 16),
    1592 => to_signed(21096, 16),
    1593 => to_signed(21057, 16),
    1594 => to_signed(21019, 16),
    1595 => to_signed(20980, 16),
    1596 => to_signed(20942, 16),
    1597 => to_signed(20903, 16),
    1598 => to_signed(20864, 16),
    1599 => to_signed(20825, 16),
    1600 => to_signed(20787, 16),
    1601 => to_signed(20748, 16),
    1602 => to_signed(20709, 16),
    1603 => to_signed(20670, 16),
    1604 => to_signed(20631, 16),
    1605 => to_signed(20592, 16),
    1606 => to_signed(20553, 16),
    1607 => to_signed(20513, 16),
    1608 => to_signed(20474, 16),
    1609 => to_signed(20435, 16),
    1610 => to_signed(20396, 16),
    1611 => to_signed(20356, 16),
    1612 => to_signed(20317, 16),
    1613 => to_signed(20277, 16),
    1614 => to_signed(20238, 16),
    1615 => to_signed(20198, 16),
    1616 => to_signed(20159, 16),
    1617 => to_signed(20119, 16),
    1618 => to_signed(20079, 16),
    1619 => to_signed(20040, 16),
    1620 => to_signed(20000, 16),
    1621 => to_signed(19960, 16),
    1622 => to_signed(19920, 16),
    1623 => to_signed(19880, 16),
    1624 => to_signed(19840, 16),
    1625 => to_signed(19800, 16),
    1626 => to_signed(19760, 16),
    1627 => to_signed(19720, 16),
    1628 => to_signed(19680, 16),
    1629 => to_signed(19640, 16),
    1630 => to_signed(19599, 16),
    1631 => to_signed(19559, 16),
    1632 => to_signed(19519, 16),
    1633 => to_signed(19478, 16),
    1634 => to_signed(19438, 16),
    1635 => to_signed(19397, 16),
    1636 => to_signed(19357, 16),
    1637 => to_signed(19316, 16),
    1638 => to_signed(19276, 16),
    1639 => to_signed(19235, 16),
    1640 => to_signed(19194, 16),
    1641 => to_signed(19154, 16),
    1642 => to_signed(19113, 16),
    1643 => to_signed(19072, 16),
    1644 => to_signed(19031, 16),
    1645 => to_signed(18990, 16),
    1646 => to_signed(18949, 16),
    1647 => to_signed(18908, 16),
    1648 => to_signed(18867, 16),
    1649 => to_signed(18826, 16),
    1650 => to_signed(18785, 16),
    1651 => to_signed(18744, 16),
    1652 => to_signed(18702, 16),
    1653 => to_signed(18661, 16),
    1654 => to_signed(18620, 16),
    1655 => to_signed(18578, 16),
    1656 => to_signed(18537, 16),
    1657 => to_signed(18495, 16),
    1658 => to_signed(18454, 16),
    1659 => to_signed(18412, 16),
    1660 => to_signed(18371, 16),
    1661 => to_signed(18329, 16),
    1662 => to_signed(18287, 16),
    1663 => to_signed(18246, 16),
    1664 => to_signed(18204, 16),
    1665 => to_signed(18162, 16),
    1666 => to_signed(18120, 16),
    1667 => to_signed(18078, 16),
    1668 => to_signed(18036, 16),
    1669 => to_signed(17994, 16),
    1670 => to_signed(17952, 16),
    1671 => to_signed(17910, 16),
    1672 => to_signed(17868, 16),
    1673 => to_signed(17826, 16),
    1674 => to_signed(17784, 16),
    1675 => to_signed(17742, 16),
    1676 => to_signed(17699, 16),
    1677 => to_signed(17657, 16),
    1678 => to_signed(17615, 16),
    1679 => to_signed(17572, 16),
    1680 => to_signed(17530, 16),
    1681 => to_signed(17487, 16),
    1682 => to_signed(17445, 16),
    1683 => to_signed(17402, 16),
    1684 => to_signed(17360, 16),
    1685 => to_signed(17317, 16),
    1686 => to_signed(17274, 16),
    1687 => to_signed(17232, 16),
    1688 => to_signed(17189, 16),
    1689 => to_signed(17146, 16),
    1690 => to_signed(17103, 16),
    1691 => to_signed(17060, 16),
    1692 => to_signed(17017, 16),
    1693 => to_signed(16974, 16),
    1694 => to_signed(16931, 16),
    1695 => to_signed(16888, 16),
    1696 => to_signed(16845, 16),
    1697 => to_signed(16802, 16),
    1698 => to_signed(16759, 16),
    1699 => to_signed(16716, 16),
    1700 => to_signed(16672, 16),
    1701 => to_signed(16629, 16),
    1702 => to_signed(16586, 16),
    1703 => to_signed(16542, 16),
    1704 => to_signed(16499, 16),
    1705 => to_signed(16455, 16),
    1706 => to_signed(16412, 16),
    1707 => to_signed(16368, 16),
    1708 => to_signed(16325, 16),
    1709 => to_signed(16281, 16),
    1710 => to_signed(16238, 16),
    1711 => to_signed(16194, 16),
    1712 => to_signed(16150, 16),
    1713 => to_signed(16107, 16),
    1714 => to_signed(16063, 16),
    1715 => to_signed(16019, 16),
    1716 => to_signed(15975, 16),
    1717 => to_signed(15931, 16),
    1718 => to_signed(15887, 16),
    1719 => to_signed(15843, 16),
    1720 => to_signed(15799, 16),
    1721 => to_signed(15755, 16),
    1722 => to_signed(15711, 16),
    1723 => to_signed(15667, 16),
    1724 => to_signed(15623, 16),
    1725 => to_signed(15579, 16),
    1726 => to_signed(15534, 16),
    1727 => to_signed(15490, 16),
    1728 => to_signed(15446, 16),
    1729 => to_signed(15401, 16),
    1730 => to_signed(15357, 16),
    1731 => to_signed(15313, 16),
    1732 => to_signed(15268, 16),
    1733 => to_signed(15224, 16),
    1734 => to_signed(15179, 16),
    1735 => to_signed(15135, 16),
    1736 => to_signed(15090, 16),
    1737 => to_signed(15045, 16),
    1738 => to_signed(15001, 16),
    1739 => to_signed(14956, 16),
    1740 => to_signed(14911, 16),
    1741 => to_signed(14866, 16),
    1742 => to_signed(14822, 16),
    1743 => to_signed(14777, 16),
    1744 => to_signed(14732, 16),
    1745 => to_signed(14687, 16),
    1746 => to_signed(14642, 16),
    1747 => to_signed(14597, 16),
    1748 => to_signed(14552, 16),
    1749 => to_signed(14507, 16),
    1750 => to_signed(14462, 16),
    1751 => to_signed(14417, 16),
    1752 => to_signed(14372, 16),
    1753 => to_signed(14326, 16),
    1754 => to_signed(14281, 16),
    1755 => to_signed(14236, 16),
    1756 => to_signed(14191, 16),
    1757 => to_signed(14145, 16),
    1758 => to_signed(14100, 16),
    1759 => to_signed(14055, 16),
    1760 => to_signed(14009, 16),
    1761 => to_signed(13964, 16),
    1762 => to_signed(13918, 16),
    1763 => to_signed(13873, 16),
    1764 => to_signed(13827, 16),
    1765 => to_signed(13782, 16),
    1766 => to_signed(13736, 16),
    1767 => to_signed(13690, 16),
    1768 => to_signed(13645, 16),
    1769 => to_signed(13599, 16),
    1770 => to_signed(13553, 16),
    1771 => to_signed(13507, 16),
    1772 => to_signed(13462, 16),
    1773 => to_signed(13416, 16),
    1774 => to_signed(13370, 16),
    1775 => to_signed(13324, 16),
    1776 => to_signed(13278, 16),
    1777 => to_signed(13232, 16),
    1778 => to_signed(13186, 16),
    1779 => to_signed(13140, 16),
    1780 => to_signed(13094, 16),
    1781 => to_signed(13048, 16),
    1782 => to_signed(13002, 16),
    1783 => to_signed(12956, 16),
    1784 => to_signed(12909, 16),
    1785 => to_signed(12863, 16),
    1786 => to_signed(12817, 16),
    1787 => to_signed(12771, 16),
    1788 => to_signed(12724, 16),
    1789 => to_signed(12678, 16),
    1790 => to_signed(12632, 16),
    1791 => to_signed(12585, 16),
    1792 => to_signed(12539, 16),
    1793 => to_signed(12492, 16),
    1794 => to_signed(12446, 16),
    1795 => to_signed(12399, 16),
    1796 => to_signed(12353, 16),
    1797 => to_signed(12306, 16),
    1798 => to_signed(12260, 16),
    1799 => to_signed(12213, 16),
    1800 => to_signed(12166, 16),
    1801 => to_signed(12120, 16),
    1802 => to_signed(12073, 16),
    1803 => to_signed(12026, 16),
    1804 => to_signed(11980, 16),
    1805 => to_signed(11933, 16),
    1806 => to_signed(11886, 16),
    1807 => to_signed(11839, 16),
    1808 => to_signed(11792, 16),
    1809 => to_signed(11745, 16),
    1810 => to_signed(11698, 16),
    1811 => to_signed(11651, 16),
    1812 => to_signed(11604, 16),
    1813 => to_signed(11557, 16),
    1814 => to_signed(11510, 16),
    1815 => to_signed(11463, 16),
    1816 => to_signed(11416, 16),
    1817 => to_signed(11369, 16),
    1818 => to_signed(11322, 16),
    1819 => to_signed(11275, 16),
    1820 => to_signed(11227, 16),
    1821 => to_signed(11180, 16),
    1822 => to_signed(11133, 16),
    1823 => to_signed(11086, 16),
    1824 => to_signed(11038, 16),
    1825 => to_signed(10991, 16),
    1826 => to_signed(10944, 16),
    1827 => to_signed(10896, 16),
    1828 => to_signed(10849, 16),
    1829 => to_signed(10801, 16),
    1830 => to_signed(10754, 16),
    1831 => to_signed(10706, 16),
    1832 => to_signed(10659, 16),
    1833 => to_signed(10611, 16),
    1834 => to_signed(10564, 16),
    1835 => to_signed(10516, 16),
    1836 => to_signed(10469, 16),
    1837 => to_signed(10421, 16),
    1838 => to_signed(10373, 16),
    1839 => to_signed(10326, 16),
    1840 => to_signed(10278, 16),
    1841 => to_signed(10230, 16),
    1842 => to_signed(10182, 16),
    1843 => to_signed(10135, 16),
    1844 => to_signed(10087, 16),
    1845 => to_signed(10039, 16),
    1846 => to_signed(9991, 16),
    1847 => to_signed(9943, 16),
    1848 => to_signed(9895, 16),
    1849 => to_signed(9847, 16),
    1850 => to_signed(9799, 16),
    1851 => to_signed(9751, 16),
    1852 => to_signed(9703, 16),
    1853 => to_signed(9655, 16),
    1854 => to_signed(9607, 16),
    1855 => to_signed(9559, 16),
    1856 => to_signed(9511, 16),
    1857 => to_signed(9463, 16),
    1858 => to_signed(9415, 16),
    1859 => to_signed(9367, 16),
    1860 => to_signed(9319, 16),
    1861 => to_signed(9270, 16),
    1862 => to_signed(9222, 16),
    1863 => to_signed(9174, 16),
    1864 => to_signed(9126, 16),
    1865 => to_signed(9077, 16),
    1866 => to_signed(9029, 16),
    1867 => to_signed(8981, 16),
    1868 => to_signed(8932, 16),
    1869 => to_signed(8884, 16),
    1870 => to_signed(8836, 16),
    1871 => to_signed(8787, 16),
    1872 => to_signed(8739, 16),
    1873 => to_signed(8690, 16),
    1874 => to_signed(8642, 16),
    1875 => to_signed(8593, 16),
    1876 => to_signed(8545, 16),
    1877 => to_signed(8496, 16),
    1878 => to_signed(8448, 16),
    1879 => to_signed(8399, 16),
    1880 => to_signed(8351, 16),
    1881 => to_signed(8302, 16),
    1882 => to_signed(8253, 16),
    1883 => to_signed(8205, 16),
    1884 => to_signed(8156, 16),
    1885 => to_signed(8107, 16),
    1886 => to_signed(8059, 16),
    1887 => to_signed(8010, 16),
    1888 => to_signed(7961, 16),
    1889 => to_signed(7912, 16),
    1890 => to_signed(7864, 16),
    1891 => to_signed(7815, 16),
    1892 => to_signed(7766, 16),
    1893 => to_signed(7717, 16),
    1894 => to_signed(7668, 16),
    1895 => to_signed(7619, 16),
    1896 => to_signed(7571, 16),
    1897 => to_signed(7522, 16),
    1898 => to_signed(7473, 16),
    1899 => to_signed(7424, 16),
    1900 => to_signed(7375, 16),
    1901 => to_signed(7326, 16),
    1902 => to_signed(7277, 16),
    1903 => to_signed(7228, 16),
    1904 => to_signed(7179, 16),
    1905 => to_signed(7130, 16),
    1906 => to_signed(7081, 16),
    1907 => to_signed(7032, 16),
    1908 => to_signed(6982, 16),
    1909 => to_signed(6933, 16),
    1910 => to_signed(6884, 16),
    1911 => to_signed(6835, 16),
    1912 => to_signed(6786, 16),
    1913 => to_signed(6737, 16),
    1914 => to_signed(6688, 16),
    1915 => to_signed(6638, 16),
    1916 => to_signed(6589, 16),
    1917 => to_signed(6540, 16),
    1918 => to_signed(6491, 16),
    1919 => to_signed(6441, 16),
    1920 => to_signed(6392, 16),
    1921 => to_signed(6343, 16),
    1922 => to_signed(6293, 16),
    1923 => to_signed(6244, 16),
    1924 => to_signed(6195, 16),
    1925 => to_signed(6145, 16),
    1926 => to_signed(6096, 16),
    1927 => to_signed(6047, 16),
    1928 => to_signed(5997, 16),
    1929 => to_signed(5948, 16),
    1930 => to_signed(5898, 16),
    1931 => to_signed(5849, 16),
    1932 => to_signed(5799, 16),
    1933 => to_signed(5750, 16),
    1934 => to_signed(5700, 16),
    1935 => to_signed(5651, 16),
    1936 => to_signed(5601, 16),
    1937 => to_signed(5552, 16),
    1938 => to_signed(5502, 16),
    1939 => to_signed(5453, 16),
    1940 => to_signed(5403, 16),
    1941 => to_signed(5354, 16),
    1942 => to_signed(5304, 16),
    1943 => to_signed(5254, 16),
    1944 => to_signed(5205, 16),
    1945 => to_signed(5155, 16),
    1946 => to_signed(5106, 16),
    1947 => to_signed(5056, 16),
    1948 => to_signed(5006, 16),
    1949 => to_signed(4957, 16),
    1950 => to_signed(4907, 16),
    1951 => to_signed(4857, 16),
    1952 => to_signed(4807, 16),
    1953 => to_signed(4758, 16),
    1954 => to_signed(4708, 16),
    1955 => to_signed(4658, 16),
    1956 => to_signed(4608, 16),
    1957 => to_signed(4559, 16),
    1958 => to_signed(4509, 16),
    1959 => to_signed(4459, 16),
    1960 => to_signed(4409, 16),
    1961 => to_signed(4359, 16),
    1962 => to_signed(4310, 16),
    1963 => to_signed(4260, 16),
    1964 => to_signed(4210, 16),
    1965 => to_signed(4160, 16),
    1966 => to_signed(4110, 16),
    1967 => to_signed(4060, 16),
    1968 => to_signed(4011, 16),
    1969 => to_signed(3961, 16),
    1970 => to_signed(3911, 16),
    1971 => to_signed(3861, 16),
    1972 => to_signed(3811, 16),
    1973 => to_signed(3761, 16),
    1974 => to_signed(3711, 16),
    1975 => to_signed(3661, 16),
    1976 => to_signed(3611, 16),
    1977 => to_signed(3561, 16),
    1978 => to_signed(3511, 16),
    1979 => to_signed(3461, 16),
    1980 => to_signed(3411, 16),
    1981 => to_signed(3361, 16),
    1982 => to_signed(3311, 16),
    1983 => to_signed(3261, 16),
    1984 => to_signed(3211, 16),
    1985 => to_signed(3161, 16),
    1986 => to_signed(3111, 16),
    1987 => to_signed(3061, 16),
    1988 => to_signed(3011, 16),
    1989 => to_signed(2961, 16),
    1990 => to_signed(2911, 16),
    1991 => to_signed(2861, 16),
    1992 => to_signed(2811, 16),
    1993 => to_signed(2761, 16),
    1994 => to_signed(2711, 16),
    1995 => to_signed(2661, 16),
    1996 => to_signed(2610, 16),
    1997 => to_signed(2560, 16),
    1998 => to_signed(2510, 16),
    1999 => to_signed(2460, 16),
    2000 => to_signed(2410, 16),
    2001 => to_signed(2360, 16),
    2002 => to_signed(2310, 16),
    2003 => to_signed(2260, 16),
    2004 => to_signed(2209, 16),
    2005 => to_signed(2159, 16),
    2006 => to_signed(2109, 16),
    2007 => to_signed(2059, 16),
    2008 => to_signed(2009, 16),
    2009 => to_signed(1959, 16),
    2010 => to_signed(1908, 16),
    2011 => to_signed(1858, 16),
    2012 => to_signed(1808, 16),
    2013 => to_signed(1758, 16),
    2014 => to_signed(1708, 16),
    2015 => to_signed(1658, 16),
    2016 => to_signed(1607, 16),
    2017 => to_signed(1557, 16),
    2018 => to_signed(1507, 16),
    2019 => to_signed(1457, 16),
    2020 => to_signed(1406, 16),
    2021 => to_signed(1356, 16),
    2022 => to_signed(1306, 16),
    2023 => to_signed(1256, 16),
    2024 => to_signed(1206, 16),
    2025 => to_signed(1155, 16),
    2026 => to_signed(1105, 16),
    2027 => to_signed(1055, 16),
    2028 => to_signed(1005, 16),
    2029 => to_signed(954, 16),
    2030 => to_signed(904, 16),
    2031 => to_signed(854, 16),
    2032 => to_signed(804, 16),
    2033 => to_signed(753, 16),
    2034 => to_signed(703, 16),
    2035 => to_signed(653, 16),
    2036 => to_signed(603, 16),
    2037 => to_signed(552, 16),
    2038 => to_signed(502, 16),
    2039 => to_signed(452, 16),
    2040 => to_signed(402, 16),
    2041 => to_signed(351, 16),
    2042 => to_signed(301, 16),
    2043 => to_signed(251, 16),
    2044 => to_signed(201, 16),
    2045 => to_signed(150, 16),
    2046 => to_signed(100, 16),
    2047 => to_signed(50, 16),
    2048 => to_signed(0, 16),
    2049 => to_signed(-50, 16),
    2050 => to_signed(-100, 16),
    2051 => to_signed(-150, 16),
    2052 => to_signed(-201, 16),
    2053 => to_signed(-251, 16),
    2054 => to_signed(-301, 16),
    2055 => to_signed(-351, 16),
    2056 => to_signed(-402, 16),
    2057 => to_signed(-452, 16),
    2058 => to_signed(-502, 16),
    2059 => to_signed(-552, 16),
    2060 => to_signed(-603, 16),
    2061 => to_signed(-653, 16),
    2062 => to_signed(-703, 16),
    2063 => to_signed(-753, 16),
    2064 => to_signed(-804, 16),
    2065 => to_signed(-854, 16),
    2066 => to_signed(-904, 16),
    2067 => to_signed(-954, 16),
    2068 => to_signed(-1005, 16),
    2069 => to_signed(-1055, 16),
    2070 => to_signed(-1105, 16),
    2071 => to_signed(-1155, 16),
    2072 => to_signed(-1206, 16),
    2073 => to_signed(-1256, 16),
    2074 => to_signed(-1306, 16),
    2075 => to_signed(-1356, 16),
    2076 => to_signed(-1406, 16),
    2077 => to_signed(-1457, 16),
    2078 => to_signed(-1507, 16),
    2079 => to_signed(-1557, 16),
    2080 => to_signed(-1607, 16),
    2081 => to_signed(-1658, 16),
    2082 => to_signed(-1708, 16),
    2083 => to_signed(-1758, 16),
    2084 => to_signed(-1808, 16),
    2085 => to_signed(-1858, 16),
    2086 => to_signed(-1908, 16),
    2087 => to_signed(-1959, 16),
    2088 => to_signed(-2009, 16),
    2089 => to_signed(-2059, 16),
    2090 => to_signed(-2109, 16),
    2091 => to_signed(-2159, 16),
    2092 => to_signed(-2209, 16),
    2093 => to_signed(-2260, 16),
    2094 => to_signed(-2310, 16),
    2095 => to_signed(-2360, 16),
    2096 => to_signed(-2410, 16),
    2097 => to_signed(-2460, 16),
    2098 => to_signed(-2510, 16),
    2099 => to_signed(-2560, 16),
    2100 => to_signed(-2610, 16),
    2101 => to_signed(-2661, 16),
    2102 => to_signed(-2711, 16),
    2103 => to_signed(-2761, 16),
    2104 => to_signed(-2811, 16),
    2105 => to_signed(-2861, 16),
    2106 => to_signed(-2911, 16),
    2107 => to_signed(-2961, 16),
    2108 => to_signed(-3011, 16),
    2109 => to_signed(-3061, 16),
    2110 => to_signed(-3111, 16),
    2111 => to_signed(-3161, 16),
    2112 => to_signed(-3211, 16),
    2113 => to_signed(-3261, 16),
    2114 => to_signed(-3311, 16),
    2115 => to_signed(-3361, 16),
    2116 => to_signed(-3411, 16),
    2117 => to_signed(-3461, 16),
    2118 => to_signed(-3511, 16),
    2119 => to_signed(-3561, 16),
    2120 => to_signed(-3611, 16),
    2121 => to_signed(-3661, 16),
    2122 => to_signed(-3711, 16),
    2123 => to_signed(-3761, 16),
    2124 => to_signed(-3811, 16),
    2125 => to_signed(-3861, 16),
    2126 => to_signed(-3911, 16),
    2127 => to_signed(-3961, 16),
    2128 => to_signed(-4011, 16),
    2129 => to_signed(-4060, 16),
    2130 => to_signed(-4110, 16),
    2131 => to_signed(-4160, 16),
    2132 => to_signed(-4210, 16),
    2133 => to_signed(-4260, 16),
    2134 => to_signed(-4310, 16),
    2135 => to_signed(-4359, 16),
    2136 => to_signed(-4409, 16),
    2137 => to_signed(-4459, 16),
    2138 => to_signed(-4509, 16),
    2139 => to_signed(-4559, 16),
    2140 => to_signed(-4608, 16),
    2141 => to_signed(-4658, 16),
    2142 => to_signed(-4708, 16),
    2143 => to_signed(-4758, 16),
    2144 => to_signed(-4807, 16),
    2145 => to_signed(-4857, 16),
    2146 => to_signed(-4907, 16),
    2147 => to_signed(-4957, 16),
    2148 => to_signed(-5006, 16),
    2149 => to_signed(-5056, 16),
    2150 => to_signed(-5106, 16),
    2151 => to_signed(-5155, 16),
    2152 => to_signed(-5205, 16),
    2153 => to_signed(-5254, 16),
    2154 => to_signed(-5304, 16),
    2155 => to_signed(-5354, 16),
    2156 => to_signed(-5403, 16),
    2157 => to_signed(-5453, 16),
    2158 => to_signed(-5502, 16),
    2159 => to_signed(-5552, 16),
    2160 => to_signed(-5601, 16),
    2161 => to_signed(-5651, 16),
    2162 => to_signed(-5700, 16),
    2163 => to_signed(-5750, 16),
    2164 => to_signed(-5799, 16),
    2165 => to_signed(-5849, 16),
    2166 => to_signed(-5898, 16),
    2167 => to_signed(-5948, 16),
    2168 => to_signed(-5997, 16),
    2169 => to_signed(-6047, 16),
    2170 => to_signed(-6096, 16),
    2171 => to_signed(-6145, 16),
    2172 => to_signed(-6195, 16),
    2173 => to_signed(-6244, 16),
    2174 => to_signed(-6293, 16),
    2175 => to_signed(-6343, 16),
    2176 => to_signed(-6392, 16),
    2177 => to_signed(-6441, 16),
    2178 => to_signed(-6491, 16),
    2179 => to_signed(-6540, 16),
    2180 => to_signed(-6589, 16),
    2181 => to_signed(-6638, 16),
    2182 => to_signed(-6688, 16),
    2183 => to_signed(-6737, 16),
    2184 => to_signed(-6786, 16),
    2185 => to_signed(-6835, 16),
    2186 => to_signed(-6884, 16),
    2187 => to_signed(-6933, 16),
    2188 => to_signed(-6982, 16),
    2189 => to_signed(-7032, 16),
    2190 => to_signed(-7081, 16),
    2191 => to_signed(-7130, 16),
    2192 => to_signed(-7179, 16),
    2193 => to_signed(-7228, 16),
    2194 => to_signed(-7277, 16),
    2195 => to_signed(-7326, 16),
    2196 => to_signed(-7375, 16),
    2197 => to_signed(-7424, 16),
    2198 => to_signed(-7473, 16),
    2199 => to_signed(-7522, 16),
    2200 => to_signed(-7571, 16),
    2201 => to_signed(-7619, 16),
    2202 => to_signed(-7668, 16),
    2203 => to_signed(-7717, 16),
    2204 => to_signed(-7766, 16),
    2205 => to_signed(-7815, 16),
    2206 => to_signed(-7864, 16),
    2207 => to_signed(-7912, 16),
    2208 => to_signed(-7961, 16),
    2209 => to_signed(-8010, 16),
    2210 => to_signed(-8059, 16),
    2211 => to_signed(-8107, 16),
    2212 => to_signed(-8156, 16),
    2213 => to_signed(-8205, 16),
    2214 => to_signed(-8253, 16),
    2215 => to_signed(-8302, 16),
    2216 => to_signed(-8351, 16),
    2217 => to_signed(-8399, 16),
    2218 => to_signed(-8448, 16),
    2219 => to_signed(-8496, 16),
    2220 => to_signed(-8545, 16),
    2221 => to_signed(-8593, 16),
    2222 => to_signed(-8642, 16),
    2223 => to_signed(-8690, 16),
    2224 => to_signed(-8739, 16),
    2225 => to_signed(-8787, 16),
    2226 => to_signed(-8836, 16),
    2227 => to_signed(-8884, 16),
    2228 => to_signed(-8932, 16),
    2229 => to_signed(-8981, 16),
    2230 => to_signed(-9029, 16),
    2231 => to_signed(-9077, 16),
    2232 => to_signed(-9126, 16),
    2233 => to_signed(-9174, 16),
    2234 => to_signed(-9222, 16),
    2235 => to_signed(-9270, 16),
    2236 => to_signed(-9319, 16),
    2237 => to_signed(-9367, 16),
    2238 => to_signed(-9415, 16),
    2239 => to_signed(-9463, 16),
    2240 => to_signed(-9511, 16),
    2241 => to_signed(-9559, 16),
    2242 => to_signed(-9607, 16),
    2243 => to_signed(-9655, 16),
    2244 => to_signed(-9703, 16),
    2245 => to_signed(-9751, 16),
    2246 => to_signed(-9799, 16),
    2247 => to_signed(-9847, 16),
    2248 => to_signed(-9895, 16),
    2249 => to_signed(-9943, 16),
    2250 => to_signed(-9991, 16),
    2251 => to_signed(-10039, 16),
    2252 => to_signed(-10087, 16),
    2253 => to_signed(-10135, 16),
    2254 => to_signed(-10182, 16),
    2255 => to_signed(-10230, 16),
    2256 => to_signed(-10278, 16),
    2257 => to_signed(-10326, 16),
    2258 => to_signed(-10373, 16),
    2259 => to_signed(-10421, 16),
    2260 => to_signed(-10469, 16),
    2261 => to_signed(-10516, 16),
    2262 => to_signed(-10564, 16),
    2263 => to_signed(-10611, 16),
    2264 => to_signed(-10659, 16),
    2265 => to_signed(-10706, 16),
    2266 => to_signed(-10754, 16),
    2267 => to_signed(-10801, 16),
    2268 => to_signed(-10849, 16),
    2269 => to_signed(-10896, 16),
    2270 => to_signed(-10944, 16),
    2271 => to_signed(-10991, 16),
    2272 => to_signed(-11038, 16),
    2273 => to_signed(-11086, 16),
    2274 => to_signed(-11133, 16),
    2275 => to_signed(-11180, 16),
    2276 => to_signed(-11227, 16),
    2277 => to_signed(-11275, 16),
    2278 => to_signed(-11322, 16),
    2279 => to_signed(-11369, 16),
    2280 => to_signed(-11416, 16),
    2281 => to_signed(-11463, 16),
    2282 => to_signed(-11510, 16),
    2283 => to_signed(-11557, 16),
    2284 => to_signed(-11604, 16),
    2285 => to_signed(-11651, 16),
    2286 => to_signed(-11698, 16),
    2287 => to_signed(-11745, 16),
    2288 => to_signed(-11792, 16),
    2289 => to_signed(-11839, 16),
    2290 => to_signed(-11886, 16),
    2291 => to_signed(-11933, 16),
    2292 => to_signed(-11980, 16),
    2293 => to_signed(-12026, 16),
    2294 => to_signed(-12073, 16),
    2295 => to_signed(-12120, 16),
    2296 => to_signed(-12166, 16),
    2297 => to_signed(-12213, 16),
    2298 => to_signed(-12260, 16),
    2299 => to_signed(-12306, 16),
    2300 => to_signed(-12353, 16),
    2301 => to_signed(-12399, 16),
    2302 => to_signed(-12446, 16),
    2303 => to_signed(-12492, 16),
    2304 => to_signed(-12539, 16),
    2305 => to_signed(-12585, 16),
    2306 => to_signed(-12632, 16),
    2307 => to_signed(-12678, 16),
    2308 => to_signed(-12724, 16),
    2309 => to_signed(-12771, 16),
    2310 => to_signed(-12817, 16),
    2311 => to_signed(-12863, 16),
    2312 => to_signed(-12909, 16),
    2313 => to_signed(-12956, 16),
    2314 => to_signed(-13002, 16),
    2315 => to_signed(-13048, 16),
    2316 => to_signed(-13094, 16),
    2317 => to_signed(-13140, 16),
    2318 => to_signed(-13186, 16),
    2319 => to_signed(-13232, 16),
    2320 => to_signed(-13278, 16),
    2321 => to_signed(-13324, 16),
    2322 => to_signed(-13370, 16),
    2323 => to_signed(-13416, 16),
    2324 => to_signed(-13462, 16),
    2325 => to_signed(-13507, 16),
    2326 => to_signed(-13553, 16),
    2327 => to_signed(-13599, 16),
    2328 => to_signed(-13645, 16),
    2329 => to_signed(-13690, 16),
    2330 => to_signed(-13736, 16),
    2331 => to_signed(-13782, 16),
    2332 => to_signed(-13827, 16),
    2333 => to_signed(-13873, 16),
    2334 => to_signed(-13918, 16),
    2335 => to_signed(-13964, 16),
    2336 => to_signed(-14009, 16),
    2337 => to_signed(-14055, 16),
    2338 => to_signed(-14100, 16),
    2339 => to_signed(-14145, 16),
    2340 => to_signed(-14191, 16),
    2341 => to_signed(-14236, 16),
    2342 => to_signed(-14281, 16),
    2343 => to_signed(-14326, 16),
    2344 => to_signed(-14372, 16),
    2345 => to_signed(-14417, 16),
    2346 => to_signed(-14462, 16),
    2347 => to_signed(-14507, 16),
    2348 => to_signed(-14552, 16),
    2349 => to_signed(-14597, 16),
    2350 => to_signed(-14642, 16),
    2351 => to_signed(-14687, 16),
    2352 => to_signed(-14732, 16),
    2353 => to_signed(-14777, 16),
    2354 => to_signed(-14822, 16),
    2355 => to_signed(-14866, 16),
    2356 => to_signed(-14911, 16),
    2357 => to_signed(-14956, 16),
    2358 => to_signed(-15001, 16),
    2359 => to_signed(-15045, 16),
    2360 => to_signed(-15090, 16),
    2361 => to_signed(-15135, 16),
    2362 => to_signed(-15179, 16),
    2363 => to_signed(-15224, 16),
    2364 => to_signed(-15268, 16),
    2365 => to_signed(-15313, 16),
    2366 => to_signed(-15357, 16),
    2367 => to_signed(-15401, 16),
    2368 => to_signed(-15446, 16),
    2369 => to_signed(-15490, 16),
    2370 => to_signed(-15534, 16),
    2371 => to_signed(-15579, 16),
    2372 => to_signed(-15623, 16),
    2373 => to_signed(-15667, 16),
    2374 => to_signed(-15711, 16),
    2375 => to_signed(-15755, 16),
    2376 => to_signed(-15799, 16),
    2377 => to_signed(-15843, 16),
    2378 => to_signed(-15887, 16),
    2379 => to_signed(-15931, 16),
    2380 => to_signed(-15975, 16),
    2381 => to_signed(-16019, 16),
    2382 => to_signed(-16063, 16),
    2383 => to_signed(-16107, 16),
    2384 => to_signed(-16150, 16),
    2385 => to_signed(-16194, 16),
    2386 => to_signed(-16238, 16),
    2387 => to_signed(-16281, 16),
    2388 => to_signed(-16325, 16),
    2389 => to_signed(-16368, 16),
    2390 => to_signed(-16412, 16),
    2391 => to_signed(-16455, 16),
    2392 => to_signed(-16499, 16),
    2393 => to_signed(-16542, 16),
    2394 => to_signed(-16586, 16),
    2395 => to_signed(-16629, 16),
    2396 => to_signed(-16672, 16),
    2397 => to_signed(-16716, 16),
    2398 => to_signed(-16759, 16),
    2399 => to_signed(-16802, 16),
    2400 => to_signed(-16845, 16),
    2401 => to_signed(-16888, 16),
    2402 => to_signed(-16931, 16),
    2403 => to_signed(-16974, 16),
    2404 => to_signed(-17017, 16),
    2405 => to_signed(-17060, 16),
    2406 => to_signed(-17103, 16),
    2407 => to_signed(-17146, 16),
    2408 => to_signed(-17189, 16),
    2409 => to_signed(-17232, 16),
    2410 => to_signed(-17274, 16),
    2411 => to_signed(-17317, 16),
    2412 => to_signed(-17360, 16),
    2413 => to_signed(-17402, 16),
    2414 => to_signed(-17445, 16),
    2415 => to_signed(-17487, 16),
    2416 => to_signed(-17530, 16),
    2417 => to_signed(-17572, 16),
    2418 => to_signed(-17615, 16),
    2419 => to_signed(-17657, 16),
    2420 => to_signed(-17699, 16),
    2421 => to_signed(-17742, 16),
    2422 => to_signed(-17784, 16),
    2423 => to_signed(-17826, 16),
    2424 => to_signed(-17868, 16),
    2425 => to_signed(-17910, 16),
    2426 => to_signed(-17952, 16),
    2427 => to_signed(-17994, 16),
    2428 => to_signed(-18036, 16),
    2429 => to_signed(-18078, 16),
    2430 => to_signed(-18120, 16),
    2431 => to_signed(-18162, 16),
    2432 => to_signed(-18204, 16),
    2433 => to_signed(-18246, 16),
    2434 => to_signed(-18287, 16),
    2435 => to_signed(-18329, 16),
    2436 => to_signed(-18371, 16),
    2437 => to_signed(-18412, 16),
    2438 => to_signed(-18454, 16),
    2439 => to_signed(-18495, 16),
    2440 => to_signed(-18537, 16),
    2441 => to_signed(-18578, 16),
    2442 => to_signed(-18620, 16),
    2443 => to_signed(-18661, 16),
    2444 => to_signed(-18702, 16),
    2445 => to_signed(-18744, 16),
    2446 => to_signed(-18785, 16),
    2447 => to_signed(-18826, 16),
    2448 => to_signed(-18867, 16),
    2449 => to_signed(-18908, 16),
    2450 => to_signed(-18949, 16),
    2451 => to_signed(-18990, 16),
    2452 => to_signed(-19031, 16),
    2453 => to_signed(-19072, 16),
    2454 => to_signed(-19113, 16),
    2455 => to_signed(-19154, 16),
    2456 => to_signed(-19194, 16),
    2457 => to_signed(-19235, 16),
    2458 => to_signed(-19276, 16),
    2459 => to_signed(-19316, 16),
    2460 => to_signed(-19357, 16),
    2461 => to_signed(-19397, 16),
    2462 => to_signed(-19438, 16),
    2463 => to_signed(-19478, 16),
    2464 => to_signed(-19519, 16),
    2465 => to_signed(-19559, 16),
    2466 => to_signed(-19599, 16),
    2467 => to_signed(-19640, 16),
    2468 => to_signed(-19680, 16),
    2469 => to_signed(-19720, 16),
    2470 => to_signed(-19760, 16),
    2471 => to_signed(-19800, 16),
    2472 => to_signed(-19840, 16),
    2473 => to_signed(-19880, 16),
    2474 => to_signed(-19920, 16),
    2475 => to_signed(-19960, 16),
    2476 => to_signed(-20000, 16),
    2477 => to_signed(-20040, 16),
    2478 => to_signed(-20079, 16),
    2479 => to_signed(-20119, 16),
    2480 => to_signed(-20159, 16),
    2481 => to_signed(-20198, 16),
    2482 => to_signed(-20238, 16),
    2483 => to_signed(-20277, 16),
    2484 => to_signed(-20317, 16),
    2485 => to_signed(-20356, 16),
    2486 => to_signed(-20396, 16),
    2487 => to_signed(-20435, 16),
    2488 => to_signed(-20474, 16),
    2489 => to_signed(-20513, 16),
    2490 => to_signed(-20553, 16),
    2491 => to_signed(-20592, 16),
    2492 => to_signed(-20631, 16),
    2493 => to_signed(-20670, 16),
    2494 => to_signed(-20709, 16),
    2495 => to_signed(-20748, 16),
    2496 => to_signed(-20787, 16),
    2497 => to_signed(-20825, 16),
    2498 => to_signed(-20864, 16),
    2499 => to_signed(-20903, 16),
    2500 => to_signed(-20942, 16),
    2501 => to_signed(-20980, 16),
    2502 => to_signed(-21019, 16),
    2503 => to_signed(-21057, 16),
    2504 => to_signed(-21096, 16),
    2505 => to_signed(-21134, 16),
    2506 => to_signed(-21173, 16),
    2507 => to_signed(-21211, 16),
    2508 => to_signed(-21249, 16),
    2509 => to_signed(-21288, 16),
    2510 => to_signed(-21326, 16),
    2511 => to_signed(-21364, 16),
    2512 => to_signed(-21402, 16),
    2513 => to_signed(-21440, 16),
    2514 => to_signed(-21478, 16),
    2515 => to_signed(-21516, 16),
    2516 => to_signed(-21554, 16),
    2517 => to_signed(-21592, 16),
    2518 => to_signed(-21629, 16),
    2519 => to_signed(-21667, 16),
    2520 => to_signed(-21705, 16),
    2521 => to_signed(-21743, 16),
    2522 => to_signed(-21780, 16),
    2523 => to_signed(-21818, 16),
    2524 => to_signed(-21855, 16),
    2525 => to_signed(-21893, 16),
    2526 => to_signed(-21930, 16),
    2527 => to_signed(-21967, 16),
    2528 => to_signed(-22004, 16),
    2529 => to_signed(-22042, 16),
    2530 => to_signed(-22079, 16),
    2531 => to_signed(-22116, 16),
    2532 => to_signed(-22153, 16),
    2533 => to_signed(-22190, 16),
    2534 => to_signed(-22227, 16),
    2535 => to_signed(-22264, 16),
    2536 => to_signed(-22301, 16),
    2537 => to_signed(-22338, 16),
    2538 => to_signed(-22374, 16),
    2539 => to_signed(-22411, 16),
    2540 => to_signed(-22448, 16),
    2541 => to_signed(-22484, 16),
    2542 => to_signed(-22521, 16),
    2543 => to_signed(-22557, 16),
    2544 => to_signed(-22594, 16),
    2545 => to_signed(-22630, 16),
    2546 => to_signed(-22666, 16),
    2547 => to_signed(-22703, 16),
    2548 => to_signed(-22739, 16),
    2549 => to_signed(-22775, 16),
    2550 => to_signed(-22811, 16),
    2551 => to_signed(-22847, 16),
    2552 => to_signed(-22883, 16),
    2553 => to_signed(-22919, 16),
    2554 => to_signed(-22955, 16),
    2555 => to_signed(-22991, 16),
    2556 => to_signed(-23027, 16),
    2557 => to_signed(-23062, 16),
    2558 => to_signed(-23098, 16),
    2559 => to_signed(-23134, 16),
    2560 => to_signed(-23169, 16),
    2561 => to_signed(-23205, 16),
    2562 => to_signed(-23240, 16),
    2563 => to_signed(-23276, 16),
    2564 => to_signed(-23311, 16),
    2565 => to_signed(-23346, 16),
    2566 => to_signed(-23382, 16),
    2567 => to_signed(-23417, 16),
    2568 => to_signed(-23452, 16),
    2569 => to_signed(-23487, 16),
    2570 => to_signed(-23522, 16),
    2571 => to_signed(-23557, 16),
    2572 => to_signed(-23592, 16),
    2573 => to_signed(-23627, 16),
    2574 => to_signed(-23661, 16),
    2575 => to_signed(-23696, 16),
    2576 => to_signed(-23731, 16),
    2577 => to_signed(-23766, 16),
    2578 => to_signed(-23800, 16),
    2579 => to_signed(-23835, 16),
    2580 => to_signed(-23869, 16),
    2581 => to_signed(-23903, 16),
    2582 => to_signed(-23938, 16),
    2583 => to_signed(-23972, 16),
    2584 => to_signed(-24006, 16),
    2585 => to_signed(-24041, 16),
    2586 => to_signed(-24075, 16),
    2587 => to_signed(-24109, 16),
    2588 => to_signed(-24143, 16),
    2589 => to_signed(-24177, 16),
    2590 => to_signed(-24211, 16),
    2591 => to_signed(-24244, 16),
    2592 => to_signed(-24278, 16),
    2593 => to_signed(-24312, 16),
    2594 => to_signed(-24346, 16),
    2595 => to_signed(-24379, 16),
    2596 => to_signed(-24413, 16),
    2597 => to_signed(-24446, 16),
    2598 => to_signed(-24480, 16),
    2599 => to_signed(-24513, 16),
    2600 => to_signed(-24546, 16),
    2601 => to_signed(-24580, 16),
    2602 => to_signed(-24613, 16),
    2603 => to_signed(-24646, 16),
    2604 => to_signed(-24679, 16),
    2605 => to_signed(-24712, 16),
    2606 => to_signed(-24745, 16),
    2607 => to_signed(-24778, 16),
    2608 => to_signed(-24811, 16),
    2609 => to_signed(-24844, 16),
    2610 => to_signed(-24877, 16),
    2611 => to_signed(-24909, 16),
    2612 => to_signed(-24942, 16),
    2613 => to_signed(-24974, 16),
    2614 => to_signed(-25007, 16),
    2615 => to_signed(-25039, 16),
    2616 => to_signed(-25072, 16),
    2617 => to_signed(-25104, 16),
    2618 => to_signed(-25136, 16),
    2619 => to_signed(-25169, 16),
    2620 => to_signed(-25201, 16),
    2621 => to_signed(-25233, 16),
    2622 => to_signed(-25265, 16),
    2623 => to_signed(-25297, 16),
    2624 => to_signed(-25329, 16),
    2625 => to_signed(-25361, 16),
    2626 => to_signed(-25392, 16),
    2627 => to_signed(-25424, 16),
    2628 => to_signed(-25456, 16),
    2629 => to_signed(-25487, 16),
    2630 => to_signed(-25519, 16),
    2631 => to_signed(-25550, 16),
    2632 => to_signed(-25582, 16),
    2633 => to_signed(-25613, 16),
    2634 => to_signed(-25645, 16),
    2635 => to_signed(-25676, 16),
    2636 => to_signed(-25707, 16),
    2637 => to_signed(-25738, 16),
    2638 => to_signed(-25769, 16),
    2639 => to_signed(-25800, 16),
    2640 => to_signed(-25831, 16),
    2641 => to_signed(-25862, 16),
    2642 => to_signed(-25893, 16),
    2643 => to_signed(-25924, 16),
    2644 => to_signed(-25954, 16),
    2645 => to_signed(-25985, 16),
    2646 => to_signed(-26016, 16),
    2647 => to_signed(-26046, 16),
    2648 => to_signed(-26077, 16),
    2649 => to_signed(-26107, 16),
    2650 => to_signed(-26137, 16),
    2651 => to_signed(-26168, 16),
    2652 => to_signed(-26198, 16),
    2653 => to_signed(-26228, 16),
    2654 => to_signed(-26258, 16),
    2655 => to_signed(-26288, 16),
    2656 => to_signed(-26318, 16),
    2657 => to_signed(-26348, 16),
    2658 => to_signed(-26378, 16),
    2659 => to_signed(-26408, 16),
    2660 => to_signed(-26437, 16),
    2661 => to_signed(-26467, 16),
    2662 => to_signed(-26497, 16),
    2663 => to_signed(-26526, 16),
    2664 => to_signed(-26556, 16),
    2665 => to_signed(-26585, 16),
    2666 => to_signed(-26615, 16),
    2667 => to_signed(-26644, 16),
    2668 => to_signed(-26673, 16),
    2669 => to_signed(-26702, 16),
    2670 => to_signed(-26731, 16),
    2671 => to_signed(-26760, 16),
    2672 => to_signed(-26789, 16),
    2673 => to_signed(-26818, 16),
    2674 => to_signed(-26847, 16),
    2675 => to_signed(-26876, 16),
    2676 => to_signed(-26905, 16),
    2677 => to_signed(-26933, 16),
    2678 => to_signed(-26962, 16),
    2679 => to_signed(-26990, 16),
    2680 => to_signed(-27019, 16),
    2681 => to_signed(-27047, 16),
    2682 => to_signed(-27076, 16),
    2683 => to_signed(-27104, 16),
    2684 => to_signed(-27132, 16),
    2685 => to_signed(-27160, 16),
    2686 => to_signed(-27188, 16),
    2687 => to_signed(-27216, 16),
    2688 => to_signed(-27244, 16),
    2689 => to_signed(-27272, 16),
    2690 => to_signed(-27300, 16),
    2691 => to_signed(-27328, 16),
    2692 => to_signed(-27355, 16),
    2693 => to_signed(-27383, 16),
    2694 => to_signed(-27411, 16),
    2695 => to_signed(-27438, 16),
    2696 => to_signed(-27466, 16),
    2697 => to_signed(-27493, 16),
    2698 => to_signed(-27520, 16),
    2699 => to_signed(-27548, 16),
    2700 => to_signed(-27575, 16),
    2701 => to_signed(-27602, 16),
    2702 => to_signed(-27629, 16),
    2703 => to_signed(-27656, 16),
    2704 => to_signed(-27683, 16),
    2705 => to_signed(-27710, 16),
    2706 => to_signed(-27736, 16),
    2707 => to_signed(-27763, 16),
    2708 => to_signed(-27790, 16),
    2709 => to_signed(-27816, 16),
    2710 => to_signed(-27843, 16),
    2711 => to_signed(-27869, 16),
    2712 => to_signed(-27896, 16),
    2713 => to_signed(-27922, 16),
    2714 => to_signed(-27948, 16),
    2715 => to_signed(-27975, 16),
    2716 => to_signed(-28001, 16),
    2717 => to_signed(-28027, 16),
    2718 => to_signed(-28053, 16),
    2719 => to_signed(-28079, 16),
    2720 => to_signed(-28105, 16),
    2721 => to_signed(-28131, 16),
    2722 => to_signed(-28156, 16),
    2723 => to_signed(-28182, 16),
    2724 => to_signed(-28208, 16),
    2725 => to_signed(-28233, 16),
    2726 => to_signed(-28259, 16),
    2727 => to_signed(-28284, 16),
    2728 => to_signed(-28309, 16),
    2729 => to_signed(-28335, 16),
    2730 => to_signed(-28360, 16),
    2731 => to_signed(-28385, 16),
    2732 => to_signed(-28410, 16),
    2733 => to_signed(-28435, 16),
    2734 => to_signed(-28460, 16),
    2735 => to_signed(-28485, 16),
    2736 => to_signed(-28510, 16),
    2737 => to_signed(-28534, 16),
    2738 => to_signed(-28559, 16),
    2739 => to_signed(-28584, 16),
    2740 => to_signed(-28608, 16),
    2741 => to_signed(-28633, 16),
    2742 => to_signed(-28657, 16),
    2743 => to_signed(-28681, 16),
    2744 => to_signed(-28706, 16),
    2745 => to_signed(-28730, 16),
    2746 => to_signed(-28754, 16),
    2747 => to_signed(-28778, 16),
    2748 => to_signed(-28802, 16),
    2749 => to_signed(-28826, 16),
    2750 => to_signed(-28850, 16),
    2751 => to_signed(-28874, 16),
    2752 => to_signed(-28897, 16),
    2753 => to_signed(-28921, 16),
    2754 => to_signed(-28945, 16),
    2755 => to_signed(-28968, 16),
    2756 => to_signed(-28992, 16),
    2757 => to_signed(-29015, 16),
    2758 => to_signed(-29038, 16),
    2759 => to_signed(-29062, 16),
    2760 => to_signed(-29085, 16),
    2761 => to_signed(-29108, 16),
    2762 => to_signed(-29131, 16),
    2763 => to_signed(-29154, 16),
    2764 => to_signed(-29177, 16),
    2765 => to_signed(-29200, 16),
    2766 => to_signed(-29222, 16),
    2767 => to_signed(-29245, 16),
    2768 => to_signed(-29268, 16),
    2769 => to_signed(-29290, 16),
    2770 => to_signed(-29313, 16),
    2771 => to_signed(-29335, 16),
    2772 => to_signed(-29358, 16),
    2773 => to_signed(-29380, 16),
    2774 => to_signed(-29402, 16),
    2775 => to_signed(-29424, 16),
    2776 => to_signed(-29446, 16),
    2777 => to_signed(-29468, 16),
    2778 => to_signed(-29490, 16),
    2779 => to_signed(-29512, 16),
    2780 => to_signed(-29534, 16),
    2781 => to_signed(-29556, 16),
    2782 => to_signed(-29577, 16),
    2783 => to_signed(-29599, 16),
    2784 => to_signed(-29621, 16),
    2785 => to_signed(-29642, 16),
    2786 => to_signed(-29663, 16),
    2787 => to_signed(-29685, 16),
    2788 => to_signed(-29706, 16),
    2789 => to_signed(-29727, 16),
    2790 => to_signed(-29748, 16),
    2791 => to_signed(-29769, 16),
    2792 => to_signed(-29790, 16),
    2793 => to_signed(-29811, 16),
    2794 => to_signed(-29832, 16),
    2795 => to_signed(-29853, 16),
    2796 => to_signed(-29873, 16),
    2797 => to_signed(-29894, 16),
    2798 => to_signed(-29915, 16),
    2799 => to_signed(-29935, 16),
    2800 => to_signed(-29955, 16),
    2801 => to_signed(-29976, 16),
    2802 => to_signed(-29996, 16),
    2803 => to_signed(-30016, 16),
    2804 => to_signed(-30036, 16),
    2805 => to_signed(-30056, 16),
    2806 => to_signed(-30076, 16),
    2807 => to_signed(-30096, 16),
    2808 => to_signed(-30116, 16),
    2809 => to_signed(-30136, 16),
    2810 => to_signed(-30156, 16),
    2811 => to_signed(-30175, 16),
    2812 => to_signed(-30195, 16),
    2813 => to_signed(-30214, 16),
    2814 => to_signed(-30234, 16),
    2815 => to_signed(-30253, 16),
    2816 => to_signed(-30272, 16),
    2817 => to_signed(-30291, 16),
    2818 => to_signed(-30311, 16),
    2819 => to_signed(-30330, 16),
    2820 => to_signed(-30349, 16),
    2821 => to_signed(-30368, 16),
    2822 => to_signed(-30386, 16),
    2823 => to_signed(-30405, 16),
    2824 => to_signed(-30424, 16),
    2825 => to_signed(-30442, 16),
    2826 => to_signed(-30461, 16),
    2827 => to_signed(-30480, 16),
    2828 => to_signed(-30498, 16),
    2829 => to_signed(-30516, 16),
    2830 => to_signed(-30535, 16),
    2831 => to_signed(-30553, 16),
    2832 => to_signed(-30571, 16),
    2833 => to_signed(-30589, 16),
    2834 => to_signed(-30607, 16),
    2835 => to_signed(-30625, 16),
    2836 => to_signed(-30643, 16),
    2837 => to_signed(-30660, 16),
    2838 => to_signed(-30678, 16),
    2839 => to_signed(-30696, 16),
    2840 => to_signed(-30713, 16),
    2841 => to_signed(-30731, 16),
    2842 => to_signed(-30748, 16),
    2843 => to_signed(-30766, 16),
    2844 => to_signed(-30783, 16),
    2845 => to_signed(-30800, 16),
    2846 => to_signed(-30817, 16),
    2847 => to_signed(-30834, 16),
    2848 => to_signed(-30851, 16),
    2849 => to_signed(-30868, 16),
    2850 => to_signed(-30885, 16),
    2851 => to_signed(-30902, 16),
    2852 => to_signed(-30918, 16),
    2853 => to_signed(-30935, 16),
    2854 => to_signed(-30951, 16),
    2855 => to_signed(-30968, 16),
    2856 => to_signed(-30984, 16),
    2857 => to_signed(-31001, 16),
    2858 => to_signed(-31017, 16),
    2859 => to_signed(-31033, 16),
    2860 => to_signed(-31049, 16),
    2861 => to_signed(-31065, 16),
    2862 => to_signed(-31081, 16),
    2863 => to_signed(-31097, 16),
    2864 => to_signed(-31113, 16),
    2865 => to_signed(-31128, 16),
    2866 => to_signed(-31144, 16),
    2867 => to_signed(-31160, 16),
    2868 => to_signed(-31175, 16),
    2869 => to_signed(-31191, 16),
    2870 => to_signed(-31206, 16),
    2871 => to_signed(-31221, 16),
    2872 => to_signed(-31236, 16),
    2873 => to_signed(-31252, 16),
    2874 => to_signed(-31267, 16),
    2875 => to_signed(-31282, 16),
    2876 => to_signed(-31297, 16),
    2877 => to_signed(-31311, 16),
    2878 => to_signed(-31326, 16),
    2879 => to_signed(-31341, 16),
    2880 => to_signed(-31356, 16),
    2881 => to_signed(-31370, 16),
    2882 => to_signed(-31385, 16),
    2883 => to_signed(-31399, 16),
    2884 => to_signed(-31413, 16),
    2885 => to_signed(-31428, 16),
    2886 => to_signed(-31442, 16),
    2887 => to_signed(-31456, 16),
    2888 => to_signed(-31470, 16),
    2889 => to_signed(-31484, 16),
    2890 => to_signed(-31498, 16),
    2891 => to_signed(-31512, 16),
    2892 => to_signed(-31525, 16),
    2893 => to_signed(-31539, 16),
    2894 => to_signed(-31553, 16),
    2895 => to_signed(-31566, 16),
    2896 => to_signed(-31580, 16),
    2897 => to_signed(-31593, 16),
    2898 => to_signed(-31606, 16),
    2899 => to_signed(-31619, 16),
    2900 => to_signed(-31633, 16),
    2901 => to_signed(-31646, 16),
    2902 => to_signed(-31659, 16),
    2903 => to_signed(-31672, 16),
    2904 => to_signed(-31684, 16),
    2905 => to_signed(-31697, 16),
    2906 => to_signed(-31710, 16),
    2907 => to_signed(-31723, 16),
    2908 => to_signed(-31735, 16),
    2909 => to_signed(-31748, 16),
    2910 => to_signed(-31760, 16),
    2911 => to_signed(-31772, 16),
    2912 => to_signed(-31785, 16),
    2913 => to_signed(-31797, 16),
    2914 => to_signed(-31809, 16),
    2915 => to_signed(-31821, 16),
    2916 => to_signed(-31833, 16),
    2917 => to_signed(-31845, 16),
    2918 => to_signed(-31856, 16),
    2919 => to_signed(-31868, 16),
    2920 => to_signed(-31880, 16),
    2921 => to_signed(-31891, 16),
    2922 => to_signed(-31903, 16),
    2923 => to_signed(-31914, 16),
    2924 => to_signed(-31926, 16),
    2925 => to_signed(-31937, 16),
    2926 => to_signed(-31948, 16),
    2927 => to_signed(-31959, 16),
    2928 => to_signed(-31970, 16),
    2929 => to_signed(-31981, 16),
    2930 => to_signed(-31992, 16),
    2931 => to_signed(-32003, 16),
    2932 => to_signed(-32014, 16),
    2933 => to_signed(-32024, 16),
    2934 => to_signed(-32035, 16),
    2935 => to_signed(-32046, 16),
    2936 => to_signed(-32056, 16),
    2937 => to_signed(-32066, 16),
    2938 => to_signed(-32077, 16),
    2939 => to_signed(-32087, 16),
    2940 => to_signed(-32097, 16),
    2941 => to_signed(-32107, 16),
    2942 => to_signed(-32117, 16),
    2943 => to_signed(-32127, 16),
    2944 => to_signed(-32137, 16),
    2945 => to_signed(-32147, 16),
    2946 => to_signed(-32156, 16),
    2947 => to_signed(-32166, 16),
    2948 => to_signed(-32176, 16),
    2949 => to_signed(-32185, 16),
    2950 => to_signed(-32194, 16),
    2951 => to_signed(-32204, 16),
    2952 => to_signed(-32213, 16),
    2953 => to_signed(-32222, 16),
    2954 => to_signed(-32231, 16),
    2955 => to_signed(-32240, 16),
    2956 => to_signed(-32249, 16),
    2957 => to_signed(-32258, 16),
    2958 => to_signed(-32267, 16),
    2959 => to_signed(-32275, 16),
    2960 => to_signed(-32284, 16),
    2961 => to_signed(-32293, 16),
    2962 => to_signed(-32301, 16),
    2963 => to_signed(-32310, 16),
    2964 => to_signed(-32318, 16),
    2965 => to_signed(-32326, 16),
    2966 => to_signed(-32334, 16),
    2967 => to_signed(-32342, 16),
    2968 => to_signed(-32350, 16),
    2969 => to_signed(-32358, 16),
    2970 => to_signed(-32366, 16),
    2971 => to_signed(-32374, 16),
    2972 => to_signed(-32382, 16),
    2973 => to_signed(-32389, 16),
    2974 => to_signed(-32397, 16),
    2975 => to_signed(-32404, 16),
    2976 => to_signed(-32412, 16),
    2977 => to_signed(-32419, 16),
    2978 => to_signed(-32426, 16),
    2979 => to_signed(-32434, 16),
    2980 => to_signed(-32441, 16),
    2981 => to_signed(-32448, 16),
    2982 => to_signed(-32455, 16),
    2983 => to_signed(-32462, 16),
    2984 => to_signed(-32468, 16),
    2985 => to_signed(-32475, 16),
    2986 => to_signed(-32482, 16),
    2987 => to_signed(-32488, 16),
    2988 => to_signed(-32495, 16),
    2989 => to_signed(-32501, 16),
    2990 => to_signed(-32508, 16),
    2991 => to_signed(-32514, 16),
    2992 => to_signed(-32520, 16),
    2993 => to_signed(-32526, 16),
    2994 => to_signed(-32532, 16),
    2995 => to_signed(-32538, 16),
    2996 => to_signed(-32544, 16),
    2997 => to_signed(-32550, 16),
    2998 => to_signed(-32556, 16),
    2999 => to_signed(-32561, 16),
    3000 => to_signed(-32567, 16),
    3001 => to_signed(-32572, 16),
    3002 => to_signed(-32578, 16),
    3003 => to_signed(-32583, 16),
    3004 => to_signed(-32588, 16),
    3005 => to_signed(-32594, 16),
    3006 => to_signed(-32599, 16),
    3007 => to_signed(-32604, 16),
    3008 => to_signed(-32609, 16),
    3009 => to_signed(-32614, 16),
    3010 => to_signed(-32618, 16),
    3011 => to_signed(-32623, 16),
    3012 => to_signed(-32628, 16),
    3013 => to_signed(-32632, 16),
    3014 => to_signed(-32637, 16),
    3015 => to_signed(-32641, 16),
    3016 => to_signed(-32646, 16),
    3017 => to_signed(-32650, 16),
    3018 => to_signed(-32654, 16),
    3019 => to_signed(-32658, 16),
    3020 => to_signed(-32662, 16),
    3021 => to_signed(-32666, 16),
    3022 => to_signed(-32670, 16),
    3023 => to_signed(-32674, 16),
    3024 => to_signed(-32678, 16),
    3025 => to_signed(-32681, 16),
    3026 => to_signed(-32685, 16),
    3027 => to_signed(-32688, 16),
    3028 => to_signed(-32692, 16),
    3029 => to_signed(-32695, 16),
    3030 => to_signed(-32699, 16),
    3031 => to_signed(-32702, 16),
    3032 => to_signed(-32705, 16),
    3033 => to_signed(-32708, 16),
    3034 => to_signed(-32711, 16),
    3035 => to_signed(-32714, 16),
    3036 => to_signed(-32717, 16),
    3037 => to_signed(-32719, 16),
    3038 => to_signed(-32722, 16),
    3039 => to_signed(-32725, 16),
    3040 => to_signed(-32727, 16),
    3041 => to_signed(-32729, 16),
    3042 => to_signed(-32732, 16),
    3043 => to_signed(-32734, 16),
    3044 => to_signed(-32736, 16),
    3045 => to_signed(-32738, 16),
    3046 => to_signed(-32740, 16),
    3047 => to_signed(-32742, 16),
    3048 => to_signed(-32744, 16),
    3049 => to_signed(-32746, 16),
    3050 => to_signed(-32748, 16),
    3051 => to_signed(-32750, 16),
    3052 => to_signed(-32751, 16),
    3053 => to_signed(-32753, 16),
    3054 => to_signed(-32754, 16),
    3055 => to_signed(-32755, 16),
    3056 => to_signed(-32757, 16),
    3057 => to_signed(-32758, 16),
    3058 => to_signed(-32759, 16),
    3059 => to_signed(-32760, 16),
    3060 => to_signed(-32761, 16),
    3061 => to_signed(-32762, 16),
    3062 => to_signed(-32763, 16),
    3063 => to_signed(-32763, 16),
    3064 => to_signed(-32764, 16),
    3065 => to_signed(-32765, 16),
    3066 => to_signed(-32765, 16),
    3067 => to_signed(-32766, 16),
    3068 => to_signed(-32766, 16),
    3069 => to_signed(-32766, 16),
    3070 => to_signed(-32766, 16),
    3071 => to_signed(-32766, 16),
    3072 => to_signed(-32767, 16),
    3073 => to_signed(-32766, 16),
    3074 => to_signed(-32766, 16),
    3075 => to_signed(-32766, 16),
    3076 => to_signed(-32766, 16),
    3077 => to_signed(-32766, 16),
    3078 => to_signed(-32765, 16),
    3079 => to_signed(-32765, 16),
    3080 => to_signed(-32764, 16),
    3081 => to_signed(-32763, 16),
    3082 => to_signed(-32763, 16),
    3083 => to_signed(-32762, 16),
    3084 => to_signed(-32761, 16),
    3085 => to_signed(-32760, 16),
    3086 => to_signed(-32759, 16),
    3087 => to_signed(-32758, 16),
    3088 => to_signed(-32757, 16),
    3089 => to_signed(-32755, 16),
    3090 => to_signed(-32754, 16),
    3091 => to_signed(-32753, 16),
    3092 => to_signed(-32751, 16),
    3093 => to_signed(-32750, 16),
    3094 => to_signed(-32748, 16),
    3095 => to_signed(-32746, 16),
    3096 => to_signed(-32744, 16),
    3097 => to_signed(-32742, 16),
    3098 => to_signed(-32740, 16),
    3099 => to_signed(-32738, 16),
    3100 => to_signed(-32736, 16),
    3101 => to_signed(-32734, 16),
    3102 => to_signed(-32732, 16),
    3103 => to_signed(-32729, 16),
    3104 => to_signed(-32727, 16),
    3105 => to_signed(-32725, 16),
    3106 => to_signed(-32722, 16),
    3107 => to_signed(-32719, 16),
    3108 => to_signed(-32717, 16),
    3109 => to_signed(-32714, 16),
    3110 => to_signed(-32711, 16),
    3111 => to_signed(-32708, 16),
    3112 => to_signed(-32705, 16),
    3113 => to_signed(-32702, 16),
    3114 => to_signed(-32699, 16),
    3115 => to_signed(-32695, 16),
    3116 => to_signed(-32692, 16),
    3117 => to_signed(-32688, 16),
    3118 => to_signed(-32685, 16),
    3119 => to_signed(-32681, 16),
    3120 => to_signed(-32678, 16),
    3121 => to_signed(-32674, 16),
    3122 => to_signed(-32670, 16),
    3123 => to_signed(-32666, 16),
    3124 => to_signed(-32662, 16),
    3125 => to_signed(-32658, 16),
    3126 => to_signed(-32654, 16),
    3127 => to_signed(-32650, 16),
    3128 => to_signed(-32646, 16),
    3129 => to_signed(-32641, 16),
    3130 => to_signed(-32637, 16),
    3131 => to_signed(-32632, 16),
    3132 => to_signed(-32628, 16),
    3133 => to_signed(-32623, 16),
    3134 => to_signed(-32618, 16),
    3135 => to_signed(-32614, 16),
    3136 => to_signed(-32609, 16),
    3137 => to_signed(-32604, 16),
    3138 => to_signed(-32599, 16),
    3139 => to_signed(-32594, 16),
    3140 => to_signed(-32588, 16),
    3141 => to_signed(-32583, 16),
    3142 => to_signed(-32578, 16),
    3143 => to_signed(-32572, 16),
    3144 => to_signed(-32567, 16),
    3145 => to_signed(-32561, 16),
    3146 => to_signed(-32556, 16),
    3147 => to_signed(-32550, 16),
    3148 => to_signed(-32544, 16),
    3149 => to_signed(-32538, 16),
    3150 => to_signed(-32532, 16),
    3151 => to_signed(-32526, 16),
    3152 => to_signed(-32520, 16),
    3153 => to_signed(-32514, 16),
    3154 => to_signed(-32508, 16),
    3155 => to_signed(-32501, 16),
    3156 => to_signed(-32495, 16),
    3157 => to_signed(-32488, 16),
    3158 => to_signed(-32482, 16),
    3159 => to_signed(-32475, 16),
    3160 => to_signed(-32468, 16),
    3161 => to_signed(-32462, 16),
    3162 => to_signed(-32455, 16),
    3163 => to_signed(-32448, 16),
    3164 => to_signed(-32441, 16),
    3165 => to_signed(-32434, 16),
    3166 => to_signed(-32426, 16),
    3167 => to_signed(-32419, 16),
    3168 => to_signed(-32412, 16),
    3169 => to_signed(-32404, 16),
    3170 => to_signed(-32397, 16),
    3171 => to_signed(-32389, 16),
    3172 => to_signed(-32382, 16),
    3173 => to_signed(-32374, 16),
    3174 => to_signed(-32366, 16),
    3175 => to_signed(-32358, 16),
    3176 => to_signed(-32350, 16),
    3177 => to_signed(-32342, 16),
    3178 => to_signed(-32334, 16),
    3179 => to_signed(-32326, 16),
    3180 => to_signed(-32318, 16),
    3181 => to_signed(-32310, 16),
    3182 => to_signed(-32301, 16),
    3183 => to_signed(-32293, 16),
    3184 => to_signed(-32284, 16),
    3185 => to_signed(-32275, 16),
    3186 => to_signed(-32267, 16),
    3187 => to_signed(-32258, 16),
    3188 => to_signed(-32249, 16),
    3189 => to_signed(-32240, 16),
    3190 => to_signed(-32231, 16),
    3191 => to_signed(-32222, 16),
    3192 => to_signed(-32213, 16),
    3193 => to_signed(-32204, 16),
    3194 => to_signed(-32194, 16),
    3195 => to_signed(-32185, 16),
    3196 => to_signed(-32176, 16),
    3197 => to_signed(-32166, 16),
    3198 => to_signed(-32156, 16),
    3199 => to_signed(-32147, 16),
    3200 => to_signed(-32137, 16),
    3201 => to_signed(-32127, 16),
    3202 => to_signed(-32117, 16),
    3203 => to_signed(-32107, 16),
    3204 => to_signed(-32097, 16),
    3205 => to_signed(-32087, 16),
    3206 => to_signed(-32077, 16),
    3207 => to_signed(-32066, 16),
    3208 => to_signed(-32056, 16),
    3209 => to_signed(-32046, 16),
    3210 => to_signed(-32035, 16),
    3211 => to_signed(-32024, 16),
    3212 => to_signed(-32014, 16),
    3213 => to_signed(-32003, 16),
    3214 => to_signed(-31992, 16),
    3215 => to_signed(-31981, 16),
    3216 => to_signed(-31970, 16),
    3217 => to_signed(-31959, 16),
    3218 => to_signed(-31948, 16),
    3219 => to_signed(-31937, 16),
    3220 => to_signed(-31926, 16),
    3221 => to_signed(-31914, 16),
    3222 => to_signed(-31903, 16),
    3223 => to_signed(-31891, 16),
    3224 => to_signed(-31880, 16),
    3225 => to_signed(-31868, 16),
    3226 => to_signed(-31856, 16),
    3227 => to_signed(-31845, 16),
    3228 => to_signed(-31833, 16),
    3229 => to_signed(-31821, 16),
    3230 => to_signed(-31809, 16),
    3231 => to_signed(-31797, 16),
    3232 => to_signed(-31785, 16),
    3233 => to_signed(-31772, 16),
    3234 => to_signed(-31760, 16),
    3235 => to_signed(-31748, 16),
    3236 => to_signed(-31735, 16),
    3237 => to_signed(-31723, 16),
    3238 => to_signed(-31710, 16),
    3239 => to_signed(-31697, 16),
    3240 => to_signed(-31684, 16),
    3241 => to_signed(-31672, 16),
    3242 => to_signed(-31659, 16),
    3243 => to_signed(-31646, 16),
    3244 => to_signed(-31633, 16),
    3245 => to_signed(-31619, 16),
    3246 => to_signed(-31606, 16),
    3247 => to_signed(-31593, 16),
    3248 => to_signed(-31580, 16),
    3249 => to_signed(-31566, 16),
    3250 => to_signed(-31553, 16),
    3251 => to_signed(-31539, 16),
    3252 => to_signed(-31525, 16),
    3253 => to_signed(-31512, 16),
    3254 => to_signed(-31498, 16),
    3255 => to_signed(-31484, 16),
    3256 => to_signed(-31470, 16),
    3257 => to_signed(-31456, 16),
    3258 => to_signed(-31442, 16),
    3259 => to_signed(-31428, 16),
    3260 => to_signed(-31413, 16),
    3261 => to_signed(-31399, 16),
    3262 => to_signed(-31385, 16),
    3263 => to_signed(-31370, 16),
    3264 => to_signed(-31356, 16),
    3265 => to_signed(-31341, 16),
    3266 => to_signed(-31326, 16),
    3267 => to_signed(-31311, 16),
    3268 => to_signed(-31297, 16),
    3269 => to_signed(-31282, 16),
    3270 => to_signed(-31267, 16),
    3271 => to_signed(-31252, 16),
    3272 => to_signed(-31236, 16),
    3273 => to_signed(-31221, 16),
    3274 => to_signed(-31206, 16),
    3275 => to_signed(-31191, 16),
    3276 => to_signed(-31175, 16),
    3277 => to_signed(-31160, 16),
    3278 => to_signed(-31144, 16),
    3279 => to_signed(-31128, 16),
    3280 => to_signed(-31113, 16),
    3281 => to_signed(-31097, 16),
    3282 => to_signed(-31081, 16),
    3283 => to_signed(-31065, 16),
    3284 => to_signed(-31049, 16),
    3285 => to_signed(-31033, 16),
    3286 => to_signed(-31017, 16),
    3287 => to_signed(-31001, 16),
    3288 => to_signed(-30984, 16),
    3289 => to_signed(-30968, 16),
    3290 => to_signed(-30951, 16),
    3291 => to_signed(-30935, 16),
    3292 => to_signed(-30918, 16),
    3293 => to_signed(-30902, 16),
    3294 => to_signed(-30885, 16),
    3295 => to_signed(-30868, 16),
    3296 => to_signed(-30851, 16),
    3297 => to_signed(-30834, 16),
    3298 => to_signed(-30817, 16),
    3299 => to_signed(-30800, 16),
    3300 => to_signed(-30783, 16),
    3301 => to_signed(-30766, 16),
    3302 => to_signed(-30748, 16),
    3303 => to_signed(-30731, 16),
    3304 => to_signed(-30713, 16),
    3305 => to_signed(-30696, 16),
    3306 => to_signed(-30678, 16),
    3307 => to_signed(-30660, 16),
    3308 => to_signed(-30643, 16),
    3309 => to_signed(-30625, 16),
    3310 => to_signed(-30607, 16),
    3311 => to_signed(-30589, 16),
    3312 => to_signed(-30571, 16),
    3313 => to_signed(-30553, 16),
    3314 => to_signed(-30535, 16),
    3315 => to_signed(-30516, 16),
    3316 => to_signed(-30498, 16),
    3317 => to_signed(-30480, 16),
    3318 => to_signed(-30461, 16),
    3319 => to_signed(-30442, 16),
    3320 => to_signed(-30424, 16),
    3321 => to_signed(-30405, 16),
    3322 => to_signed(-30386, 16),
    3323 => to_signed(-30368, 16),
    3324 => to_signed(-30349, 16),
    3325 => to_signed(-30330, 16),
    3326 => to_signed(-30311, 16),
    3327 => to_signed(-30291, 16),
    3328 => to_signed(-30272, 16),
    3329 => to_signed(-30253, 16),
    3330 => to_signed(-30234, 16),
    3331 => to_signed(-30214, 16),
    3332 => to_signed(-30195, 16),
    3333 => to_signed(-30175, 16),
    3334 => to_signed(-30156, 16),
    3335 => to_signed(-30136, 16),
    3336 => to_signed(-30116, 16),
    3337 => to_signed(-30096, 16),
    3338 => to_signed(-30076, 16),
    3339 => to_signed(-30056, 16),
    3340 => to_signed(-30036, 16),
    3341 => to_signed(-30016, 16),
    3342 => to_signed(-29996, 16),
    3343 => to_signed(-29976, 16),
    3344 => to_signed(-29955, 16),
    3345 => to_signed(-29935, 16),
    3346 => to_signed(-29915, 16),
    3347 => to_signed(-29894, 16),
    3348 => to_signed(-29873, 16),
    3349 => to_signed(-29853, 16),
    3350 => to_signed(-29832, 16),
    3351 => to_signed(-29811, 16),
    3352 => to_signed(-29790, 16),
    3353 => to_signed(-29769, 16),
    3354 => to_signed(-29748, 16),
    3355 => to_signed(-29727, 16),
    3356 => to_signed(-29706, 16),
    3357 => to_signed(-29685, 16),
    3358 => to_signed(-29663, 16),
    3359 => to_signed(-29642, 16),
    3360 => to_signed(-29621, 16),
    3361 => to_signed(-29599, 16),
    3362 => to_signed(-29577, 16),
    3363 => to_signed(-29556, 16),
    3364 => to_signed(-29534, 16),
    3365 => to_signed(-29512, 16),
    3366 => to_signed(-29490, 16),
    3367 => to_signed(-29468, 16),
    3368 => to_signed(-29446, 16),
    3369 => to_signed(-29424, 16),
    3370 => to_signed(-29402, 16),
    3371 => to_signed(-29380, 16),
    3372 => to_signed(-29358, 16),
    3373 => to_signed(-29335, 16),
    3374 => to_signed(-29313, 16),
    3375 => to_signed(-29290, 16),
    3376 => to_signed(-29268, 16),
    3377 => to_signed(-29245, 16),
    3378 => to_signed(-29222, 16),
    3379 => to_signed(-29200, 16),
    3380 => to_signed(-29177, 16),
    3381 => to_signed(-29154, 16),
    3382 => to_signed(-29131, 16),
    3383 => to_signed(-29108, 16),
    3384 => to_signed(-29085, 16),
    3385 => to_signed(-29062, 16),
    3386 => to_signed(-29038, 16),
    3387 => to_signed(-29015, 16),
    3388 => to_signed(-28992, 16),
    3389 => to_signed(-28968, 16),
    3390 => to_signed(-28945, 16),
    3391 => to_signed(-28921, 16),
    3392 => to_signed(-28897, 16),
    3393 => to_signed(-28874, 16),
    3394 => to_signed(-28850, 16),
    3395 => to_signed(-28826, 16),
    3396 => to_signed(-28802, 16),
    3397 => to_signed(-28778, 16),
    3398 => to_signed(-28754, 16),
    3399 => to_signed(-28730, 16),
    3400 => to_signed(-28706, 16),
    3401 => to_signed(-28681, 16),
    3402 => to_signed(-28657, 16),
    3403 => to_signed(-28633, 16),
    3404 => to_signed(-28608, 16),
    3405 => to_signed(-28584, 16),
    3406 => to_signed(-28559, 16),
    3407 => to_signed(-28534, 16),
    3408 => to_signed(-28510, 16),
    3409 => to_signed(-28485, 16),
    3410 => to_signed(-28460, 16),
    3411 => to_signed(-28435, 16),
    3412 => to_signed(-28410, 16),
    3413 => to_signed(-28385, 16),
    3414 => to_signed(-28360, 16),
    3415 => to_signed(-28335, 16),
    3416 => to_signed(-28309, 16),
    3417 => to_signed(-28284, 16),
    3418 => to_signed(-28259, 16),
    3419 => to_signed(-28233, 16),
    3420 => to_signed(-28208, 16),
    3421 => to_signed(-28182, 16),
    3422 => to_signed(-28156, 16),
    3423 => to_signed(-28131, 16),
    3424 => to_signed(-28105, 16),
    3425 => to_signed(-28079, 16),
    3426 => to_signed(-28053, 16),
    3427 => to_signed(-28027, 16),
    3428 => to_signed(-28001, 16),
    3429 => to_signed(-27975, 16),
    3430 => to_signed(-27948, 16),
    3431 => to_signed(-27922, 16),
    3432 => to_signed(-27896, 16),
    3433 => to_signed(-27869, 16),
    3434 => to_signed(-27843, 16),
    3435 => to_signed(-27816, 16),
    3436 => to_signed(-27790, 16),
    3437 => to_signed(-27763, 16),
    3438 => to_signed(-27736, 16),
    3439 => to_signed(-27710, 16),
    3440 => to_signed(-27683, 16),
    3441 => to_signed(-27656, 16),
    3442 => to_signed(-27629, 16),
    3443 => to_signed(-27602, 16),
    3444 => to_signed(-27575, 16),
    3445 => to_signed(-27548, 16),
    3446 => to_signed(-27520, 16),
    3447 => to_signed(-27493, 16),
    3448 => to_signed(-27466, 16),
    3449 => to_signed(-27438, 16),
    3450 => to_signed(-27411, 16),
    3451 => to_signed(-27383, 16),
    3452 => to_signed(-27355, 16),
    3453 => to_signed(-27328, 16),
    3454 => to_signed(-27300, 16),
    3455 => to_signed(-27272, 16),
    3456 => to_signed(-27244, 16),
    3457 => to_signed(-27216, 16),
    3458 => to_signed(-27188, 16),
    3459 => to_signed(-27160, 16),
    3460 => to_signed(-27132, 16),
    3461 => to_signed(-27104, 16),
    3462 => to_signed(-27076, 16),
    3463 => to_signed(-27047, 16),
    3464 => to_signed(-27019, 16),
    3465 => to_signed(-26990, 16),
    3466 => to_signed(-26962, 16),
    3467 => to_signed(-26933, 16),
    3468 => to_signed(-26905, 16),
    3469 => to_signed(-26876, 16),
    3470 => to_signed(-26847, 16),
    3471 => to_signed(-26818, 16),
    3472 => to_signed(-26789, 16),
    3473 => to_signed(-26760, 16),
    3474 => to_signed(-26731, 16),
    3475 => to_signed(-26702, 16),
    3476 => to_signed(-26673, 16),
    3477 => to_signed(-26644, 16),
    3478 => to_signed(-26615, 16),
    3479 => to_signed(-26585, 16),
    3480 => to_signed(-26556, 16),
    3481 => to_signed(-26526, 16),
    3482 => to_signed(-26497, 16),
    3483 => to_signed(-26467, 16),
    3484 => to_signed(-26437, 16),
    3485 => to_signed(-26408, 16),
    3486 => to_signed(-26378, 16),
    3487 => to_signed(-26348, 16),
    3488 => to_signed(-26318, 16),
    3489 => to_signed(-26288, 16),
    3490 => to_signed(-26258, 16),
    3491 => to_signed(-26228, 16),
    3492 => to_signed(-26198, 16),
    3493 => to_signed(-26168, 16),
    3494 => to_signed(-26137, 16),
    3495 => to_signed(-26107, 16),
    3496 => to_signed(-26077, 16),
    3497 => to_signed(-26046, 16),
    3498 => to_signed(-26016, 16),
    3499 => to_signed(-25985, 16),
    3500 => to_signed(-25954, 16),
    3501 => to_signed(-25924, 16),
    3502 => to_signed(-25893, 16),
    3503 => to_signed(-25862, 16),
    3504 => to_signed(-25831, 16),
    3505 => to_signed(-25800, 16),
    3506 => to_signed(-25769, 16),
    3507 => to_signed(-25738, 16),
    3508 => to_signed(-25707, 16),
    3509 => to_signed(-25676, 16),
    3510 => to_signed(-25645, 16),
    3511 => to_signed(-25613, 16),
    3512 => to_signed(-25582, 16),
    3513 => to_signed(-25550, 16),
    3514 => to_signed(-25519, 16),
    3515 => to_signed(-25487, 16),
    3516 => to_signed(-25456, 16),
    3517 => to_signed(-25424, 16),
    3518 => to_signed(-25392, 16),
    3519 => to_signed(-25361, 16),
    3520 => to_signed(-25329, 16),
    3521 => to_signed(-25297, 16),
    3522 => to_signed(-25265, 16),
    3523 => to_signed(-25233, 16),
    3524 => to_signed(-25201, 16),
    3525 => to_signed(-25169, 16),
    3526 => to_signed(-25136, 16),
    3527 => to_signed(-25104, 16),
    3528 => to_signed(-25072, 16),
    3529 => to_signed(-25039, 16),
    3530 => to_signed(-25007, 16),
    3531 => to_signed(-24974, 16),
    3532 => to_signed(-24942, 16),
    3533 => to_signed(-24909, 16),
    3534 => to_signed(-24877, 16),
    3535 => to_signed(-24844, 16),
    3536 => to_signed(-24811, 16),
    3537 => to_signed(-24778, 16),
    3538 => to_signed(-24745, 16),
    3539 => to_signed(-24712, 16),
    3540 => to_signed(-24679, 16),
    3541 => to_signed(-24646, 16),
    3542 => to_signed(-24613, 16),
    3543 => to_signed(-24580, 16),
    3544 => to_signed(-24546, 16),
    3545 => to_signed(-24513, 16),
    3546 => to_signed(-24480, 16),
    3547 => to_signed(-24446, 16),
    3548 => to_signed(-24413, 16),
    3549 => to_signed(-24379, 16),
    3550 => to_signed(-24346, 16),
    3551 => to_signed(-24312, 16),
    3552 => to_signed(-24278, 16),
    3553 => to_signed(-24244, 16),
    3554 => to_signed(-24211, 16),
    3555 => to_signed(-24177, 16),
    3556 => to_signed(-24143, 16),
    3557 => to_signed(-24109, 16),
    3558 => to_signed(-24075, 16),
    3559 => to_signed(-24041, 16),
    3560 => to_signed(-24006, 16),
    3561 => to_signed(-23972, 16),
    3562 => to_signed(-23938, 16),
    3563 => to_signed(-23903, 16),
    3564 => to_signed(-23869, 16),
    3565 => to_signed(-23835, 16),
    3566 => to_signed(-23800, 16),
    3567 => to_signed(-23766, 16),
    3568 => to_signed(-23731, 16),
    3569 => to_signed(-23696, 16),
    3570 => to_signed(-23661, 16),
    3571 => to_signed(-23627, 16),
    3572 => to_signed(-23592, 16),
    3573 => to_signed(-23557, 16),
    3574 => to_signed(-23522, 16),
    3575 => to_signed(-23487, 16),
    3576 => to_signed(-23452, 16),
    3577 => to_signed(-23417, 16),
    3578 => to_signed(-23382, 16),
    3579 => to_signed(-23346, 16),
    3580 => to_signed(-23311, 16),
    3581 => to_signed(-23276, 16),
    3582 => to_signed(-23240, 16),
    3583 => to_signed(-23205, 16),
    3584 => to_signed(-23169, 16),
    3585 => to_signed(-23134, 16),
    3586 => to_signed(-23098, 16),
    3587 => to_signed(-23062, 16),
    3588 => to_signed(-23027, 16),
    3589 => to_signed(-22991, 16),
    3590 => to_signed(-22955, 16),
    3591 => to_signed(-22919, 16),
    3592 => to_signed(-22883, 16),
    3593 => to_signed(-22847, 16),
    3594 => to_signed(-22811, 16),
    3595 => to_signed(-22775, 16),
    3596 => to_signed(-22739, 16),
    3597 => to_signed(-22703, 16),
    3598 => to_signed(-22666, 16),
    3599 => to_signed(-22630, 16),
    3600 => to_signed(-22594, 16),
    3601 => to_signed(-22557, 16),
    3602 => to_signed(-22521, 16),
    3603 => to_signed(-22484, 16),
    3604 => to_signed(-22448, 16),
    3605 => to_signed(-22411, 16),
    3606 => to_signed(-22374, 16),
    3607 => to_signed(-22338, 16),
    3608 => to_signed(-22301, 16),
    3609 => to_signed(-22264, 16),
    3610 => to_signed(-22227, 16),
    3611 => to_signed(-22190, 16),
    3612 => to_signed(-22153, 16),
    3613 => to_signed(-22116, 16),
    3614 => to_signed(-22079, 16),
    3615 => to_signed(-22042, 16),
    3616 => to_signed(-22004, 16),
    3617 => to_signed(-21967, 16),
    3618 => to_signed(-21930, 16),
    3619 => to_signed(-21893, 16),
    3620 => to_signed(-21855, 16),
    3621 => to_signed(-21818, 16),
    3622 => to_signed(-21780, 16),
    3623 => to_signed(-21743, 16),
    3624 => to_signed(-21705, 16),
    3625 => to_signed(-21667, 16),
    3626 => to_signed(-21629, 16),
    3627 => to_signed(-21592, 16),
    3628 => to_signed(-21554, 16),
    3629 => to_signed(-21516, 16),
    3630 => to_signed(-21478, 16),
    3631 => to_signed(-21440, 16),
    3632 => to_signed(-21402, 16),
    3633 => to_signed(-21364, 16),
    3634 => to_signed(-21326, 16),
    3635 => to_signed(-21288, 16),
    3636 => to_signed(-21249, 16),
    3637 => to_signed(-21211, 16),
    3638 => to_signed(-21173, 16),
    3639 => to_signed(-21134, 16),
    3640 => to_signed(-21096, 16),
    3641 => to_signed(-21057, 16),
    3642 => to_signed(-21019, 16),
    3643 => to_signed(-20980, 16),
    3644 => to_signed(-20942, 16),
    3645 => to_signed(-20903, 16),
    3646 => to_signed(-20864, 16),
    3647 => to_signed(-20825, 16),
    3648 => to_signed(-20787, 16),
    3649 => to_signed(-20748, 16),
    3650 => to_signed(-20709, 16),
    3651 => to_signed(-20670, 16),
    3652 => to_signed(-20631, 16),
    3653 => to_signed(-20592, 16),
    3654 => to_signed(-20553, 16),
    3655 => to_signed(-20513, 16),
    3656 => to_signed(-20474, 16),
    3657 => to_signed(-20435, 16),
    3658 => to_signed(-20396, 16),
    3659 => to_signed(-20356, 16),
    3660 => to_signed(-20317, 16),
    3661 => to_signed(-20277, 16),
    3662 => to_signed(-20238, 16),
    3663 => to_signed(-20198, 16),
    3664 => to_signed(-20159, 16),
    3665 => to_signed(-20119, 16),
    3666 => to_signed(-20079, 16),
    3667 => to_signed(-20040, 16),
    3668 => to_signed(-20000, 16),
    3669 => to_signed(-19960, 16),
    3670 => to_signed(-19920, 16),
    3671 => to_signed(-19880, 16),
    3672 => to_signed(-19840, 16),
    3673 => to_signed(-19800, 16),
    3674 => to_signed(-19760, 16),
    3675 => to_signed(-19720, 16),
    3676 => to_signed(-19680, 16),
    3677 => to_signed(-19640, 16),
    3678 => to_signed(-19599, 16),
    3679 => to_signed(-19559, 16),
    3680 => to_signed(-19519, 16),
    3681 => to_signed(-19478, 16),
    3682 => to_signed(-19438, 16),
    3683 => to_signed(-19397, 16),
    3684 => to_signed(-19357, 16),
    3685 => to_signed(-19316, 16),
    3686 => to_signed(-19276, 16),
    3687 => to_signed(-19235, 16),
    3688 => to_signed(-19194, 16),
    3689 => to_signed(-19154, 16),
    3690 => to_signed(-19113, 16),
    3691 => to_signed(-19072, 16),
    3692 => to_signed(-19031, 16),
    3693 => to_signed(-18990, 16),
    3694 => to_signed(-18949, 16),
    3695 => to_signed(-18908, 16),
    3696 => to_signed(-18867, 16),
    3697 => to_signed(-18826, 16),
    3698 => to_signed(-18785, 16),
    3699 => to_signed(-18744, 16),
    3700 => to_signed(-18702, 16),
    3701 => to_signed(-18661, 16),
    3702 => to_signed(-18620, 16),
    3703 => to_signed(-18578, 16),
    3704 => to_signed(-18537, 16),
    3705 => to_signed(-18495, 16),
    3706 => to_signed(-18454, 16),
    3707 => to_signed(-18412, 16),
    3708 => to_signed(-18371, 16),
    3709 => to_signed(-18329, 16),
    3710 => to_signed(-18287, 16),
    3711 => to_signed(-18246, 16),
    3712 => to_signed(-18204, 16),
    3713 => to_signed(-18162, 16),
    3714 => to_signed(-18120, 16),
    3715 => to_signed(-18078, 16),
    3716 => to_signed(-18036, 16),
    3717 => to_signed(-17994, 16),
    3718 => to_signed(-17952, 16),
    3719 => to_signed(-17910, 16),
    3720 => to_signed(-17868, 16),
    3721 => to_signed(-17826, 16),
    3722 => to_signed(-17784, 16),
    3723 => to_signed(-17742, 16),
    3724 => to_signed(-17699, 16),
    3725 => to_signed(-17657, 16),
    3726 => to_signed(-17615, 16),
    3727 => to_signed(-17572, 16),
    3728 => to_signed(-17530, 16),
    3729 => to_signed(-17487, 16),
    3730 => to_signed(-17445, 16),
    3731 => to_signed(-17402, 16),
    3732 => to_signed(-17360, 16),
    3733 => to_signed(-17317, 16),
    3734 => to_signed(-17274, 16),
    3735 => to_signed(-17232, 16),
    3736 => to_signed(-17189, 16),
    3737 => to_signed(-17146, 16),
    3738 => to_signed(-17103, 16),
    3739 => to_signed(-17060, 16),
    3740 => to_signed(-17017, 16),
    3741 => to_signed(-16974, 16),
    3742 => to_signed(-16931, 16),
    3743 => to_signed(-16888, 16),
    3744 => to_signed(-16845, 16),
    3745 => to_signed(-16802, 16),
    3746 => to_signed(-16759, 16),
    3747 => to_signed(-16716, 16),
    3748 => to_signed(-16672, 16),
    3749 => to_signed(-16629, 16),
    3750 => to_signed(-16586, 16),
    3751 => to_signed(-16542, 16),
    3752 => to_signed(-16499, 16),
    3753 => to_signed(-16455, 16),
    3754 => to_signed(-16412, 16),
    3755 => to_signed(-16368, 16),
    3756 => to_signed(-16325, 16),
    3757 => to_signed(-16281, 16),
    3758 => to_signed(-16238, 16),
    3759 => to_signed(-16194, 16),
    3760 => to_signed(-16150, 16),
    3761 => to_signed(-16107, 16),
    3762 => to_signed(-16063, 16),
    3763 => to_signed(-16019, 16),
    3764 => to_signed(-15975, 16),
    3765 => to_signed(-15931, 16),
    3766 => to_signed(-15887, 16),
    3767 => to_signed(-15843, 16),
    3768 => to_signed(-15799, 16),
    3769 => to_signed(-15755, 16),
    3770 => to_signed(-15711, 16),
    3771 => to_signed(-15667, 16),
    3772 => to_signed(-15623, 16),
    3773 => to_signed(-15579, 16),
    3774 => to_signed(-15534, 16),
    3775 => to_signed(-15490, 16),
    3776 => to_signed(-15446, 16),
    3777 => to_signed(-15401, 16),
    3778 => to_signed(-15357, 16),
    3779 => to_signed(-15313, 16),
    3780 => to_signed(-15268, 16),
    3781 => to_signed(-15224, 16),
    3782 => to_signed(-15179, 16),
    3783 => to_signed(-15135, 16),
    3784 => to_signed(-15090, 16),
    3785 => to_signed(-15045, 16),
    3786 => to_signed(-15001, 16),
    3787 => to_signed(-14956, 16),
    3788 => to_signed(-14911, 16),
    3789 => to_signed(-14866, 16),
    3790 => to_signed(-14822, 16),
    3791 => to_signed(-14777, 16),
    3792 => to_signed(-14732, 16),
    3793 => to_signed(-14687, 16),
    3794 => to_signed(-14642, 16),
    3795 => to_signed(-14597, 16),
    3796 => to_signed(-14552, 16),
    3797 => to_signed(-14507, 16),
    3798 => to_signed(-14462, 16),
    3799 => to_signed(-14417, 16),
    3800 => to_signed(-14372, 16),
    3801 => to_signed(-14326, 16),
    3802 => to_signed(-14281, 16),
    3803 => to_signed(-14236, 16),
    3804 => to_signed(-14191, 16),
    3805 => to_signed(-14145, 16),
    3806 => to_signed(-14100, 16),
    3807 => to_signed(-14055, 16),
    3808 => to_signed(-14009, 16),
    3809 => to_signed(-13964, 16),
    3810 => to_signed(-13918, 16),
    3811 => to_signed(-13873, 16),
    3812 => to_signed(-13827, 16),
    3813 => to_signed(-13782, 16),
    3814 => to_signed(-13736, 16),
    3815 => to_signed(-13690, 16),
    3816 => to_signed(-13645, 16),
    3817 => to_signed(-13599, 16),
    3818 => to_signed(-13553, 16),
    3819 => to_signed(-13507, 16),
    3820 => to_signed(-13462, 16),
    3821 => to_signed(-13416, 16),
    3822 => to_signed(-13370, 16),
    3823 => to_signed(-13324, 16),
    3824 => to_signed(-13278, 16),
    3825 => to_signed(-13232, 16),
    3826 => to_signed(-13186, 16),
    3827 => to_signed(-13140, 16),
    3828 => to_signed(-13094, 16),
    3829 => to_signed(-13048, 16),
    3830 => to_signed(-13002, 16),
    3831 => to_signed(-12956, 16),
    3832 => to_signed(-12909, 16),
    3833 => to_signed(-12863, 16),
    3834 => to_signed(-12817, 16),
    3835 => to_signed(-12771, 16),
    3836 => to_signed(-12724, 16),
    3837 => to_signed(-12678, 16),
    3838 => to_signed(-12632, 16),
    3839 => to_signed(-12585, 16),
    3840 => to_signed(-12539, 16),
    3841 => to_signed(-12492, 16),
    3842 => to_signed(-12446, 16),
    3843 => to_signed(-12399, 16),
    3844 => to_signed(-12353, 16),
    3845 => to_signed(-12306, 16),
    3846 => to_signed(-12260, 16),
    3847 => to_signed(-12213, 16),
    3848 => to_signed(-12166, 16),
    3849 => to_signed(-12120, 16),
    3850 => to_signed(-12073, 16),
    3851 => to_signed(-12026, 16),
    3852 => to_signed(-11980, 16),
    3853 => to_signed(-11933, 16),
    3854 => to_signed(-11886, 16),
    3855 => to_signed(-11839, 16),
    3856 => to_signed(-11792, 16),
    3857 => to_signed(-11745, 16),
    3858 => to_signed(-11698, 16),
    3859 => to_signed(-11651, 16),
    3860 => to_signed(-11604, 16),
    3861 => to_signed(-11557, 16),
    3862 => to_signed(-11510, 16),
    3863 => to_signed(-11463, 16),
    3864 => to_signed(-11416, 16),
    3865 => to_signed(-11369, 16),
    3866 => to_signed(-11322, 16),
    3867 => to_signed(-11275, 16),
    3868 => to_signed(-11227, 16),
    3869 => to_signed(-11180, 16),
    3870 => to_signed(-11133, 16),
    3871 => to_signed(-11086, 16),
    3872 => to_signed(-11038, 16),
    3873 => to_signed(-10991, 16),
    3874 => to_signed(-10944, 16),
    3875 => to_signed(-10896, 16),
    3876 => to_signed(-10849, 16),
    3877 => to_signed(-10801, 16),
    3878 => to_signed(-10754, 16),
    3879 => to_signed(-10706, 16),
    3880 => to_signed(-10659, 16),
    3881 => to_signed(-10611, 16),
    3882 => to_signed(-10564, 16),
    3883 => to_signed(-10516, 16),
    3884 => to_signed(-10469, 16),
    3885 => to_signed(-10421, 16),
    3886 => to_signed(-10373, 16),
    3887 => to_signed(-10326, 16),
    3888 => to_signed(-10278, 16),
    3889 => to_signed(-10230, 16),
    3890 => to_signed(-10182, 16),
    3891 => to_signed(-10135, 16),
    3892 => to_signed(-10087, 16),
    3893 => to_signed(-10039, 16),
    3894 => to_signed(-9991, 16),
    3895 => to_signed(-9943, 16),
    3896 => to_signed(-9895, 16),
    3897 => to_signed(-9847, 16),
    3898 => to_signed(-9799, 16),
    3899 => to_signed(-9751, 16),
    3900 => to_signed(-9703, 16),
    3901 => to_signed(-9655, 16),
    3902 => to_signed(-9607, 16),
    3903 => to_signed(-9559, 16),
    3904 => to_signed(-9511, 16),
    3905 => to_signed(-9463, 16),
    3906 => to_signed(-9415, 16),
    3907 => to_signed(-9367, 16),
    3908 => to_signed(-9319, 16),
    3909 => to_signed(-9270, 16),
    3910 => to_signed(-9222, 16),
    3911 => to_signed(-9174, 16),
    3912 => to_signed(-9126, 16),
    3913 => to_signed(-9077, 16),
    3914 => to_signed(-9029, 16),
    3915 => to_signed(-8981, 16),
    3916 => to_signed(-8932, 16),
    3917 => to_signed(-8884, 16),
    3918 => to_signed(-8836, 16),
    3919 => to_signed(-8787, 16),
    3920 => to_signed(-8739, 16),
    3921 => to_signed(-8690, 16),
    3922 => to_signed(-8642, 16),
    3923 => to_signed(-8593, 16),
    3924 => to_signed(-8545, 16),
    3925 => to_signed(-8496, 16),
    3926 => to_signed(-8448, 16),
    3927 => to_signed(-8399, 16),
    3928 => to_signed(-8351, 16),
    3929 => to_signed(-8302, 16),
    3930 => to_signed(-8253, 16),
    3931 => to_signed(-8205, 16),
    3932 => to_signed(-8156, 16),
    3933 => to_signed(-8107, 16),
    3934 => to_signed(-8059, 16),
    3935 => to_signed(-8010, 16),
    3936 => to_signed(-7961, 16),
    3937 => to_signed(-7912, 16),
    3938 => to_signed(-7864, 16),
    3939 => to_signed(-7815, 16),
    3940 => to_signed(-7766, 16),
    3941 => to_signed(-7717, 16),
    3942 => to_signed(-7668, 16),
    3943 => to_signed(-7619, 16),
    3944 => to_signed(-7571, 16),
    3945 => to_signed(-7522, 16),
    3946 => to_signed(-7473, 16),
    3947 => to_signed(-7424, 16),
    3948 => to_signed(-7375, 16),
    3949 => to_signed(-7326, 16),
    3950 => to_signed(-7277, 16),
    3951 => to_signed(-7228, 16),
    3952 => to_signed(-7179, 16),
    3953 => to_signed(-7130, 16),
    3954 => to_signed(-7081, 16),
    3955 => to_signed(-7032, 16),
    3956 => to_signed(-6982, 16),
    3957 => to_signed(-6933, 16),
    3958 => to_signed(-6884, 16),
    3959 => to_signed(-6835, 16),
    3960 => to_signed(-6786, 16),
    3961 => to_signed(-6737, 16),
    3962 => to_signed(-6688, 16),
    3963 => to_signed(-6638, 16),
    3964 => to_signed(-6589, 16),
    3965 => to_signed(-6540, 16),
    3966 => to_signed(-6491, 16),
    3967 => to_signed(-6441, 16),
    3968 => to_signed(-6392, 16),
    3969 => to_signed(-6343, 16),
    3970 => to_signed(-6293, 16),
    3971 => to_signed(-6244, 16),
    3972 => to_signed(-6195, 16),
    3973 => to_signed(-6145, 16),
    3974 => to_signed(-6096, 16),
    3975 => to_signed(-6047, 16),
    3976 => to_signed(-5997, 16),
    3977 => to_signed(-5948, 16),
    3978 => to_signed(-5898, 16),
    3979 => to_signed(-5849, 16),
    3980 => to_signed(-5799, 16),
    3981 => to_signed(-5750, 16),
    3982 => to_signed(-5700, 16),
    3983 => to_signed(-5651, 16),
    3984 => to_signed(-5601, 16),
    3985 => to_signed(-5552, 16),
    3986 => to_signed(-5502, 16),
    3987 => to_signed(-5453, 16),
    3988 => to_signed(-5403, 16),
    3989 => to_signed(-5354, 16),
    3990 => to_signed(-5304, 16),
    3991 => to_signed(-5254, 16),
    3992 => to_signed(-5205, 16),
    3993 => to_signed(-5155, 16),
    3994 => to_signed(-5106, 16),
    3995 => to_signed(-5056, 16),
    3996 => to_signed(-5006, 16),
    3997 => to_signed(-4957, 16),
    3998 => to_signed(-4907, 16),
    3999 => to_signed(-4857, 16),
    4000 => to_signed(-4807, 16),
    4001 => to_signed(-4758, 16),
    4002 => to_signed(-4708, 16),
    4003 => to_signed(-4658, 16),
    4004 => to_signed(-4608, 16),
    4005 => to_signed(-4559, 16),
    4006 => to_signed(-4509, 16),
    4007 => to_signed(-4459, 16),
    4008 => to_signed(-4409, 16),
    4009 => to_signed(-4359, 16),
    4010 => to_signed(-4310, 16),
    4011 => to_signed(-4260, 16),
    4012 => to_signed(-4210, 16),
    4013 => to_signed(-4160, 16),
    4014 => to_signed(-4110, 16),
    4015 => to_signed(-4060, 16),
    4016 => to_signed(-4011, 16),
    4017 => to_signed(-3961, 16),
    4018 => to_signed(-3911, 16),
    4019 => to_signed(-3861, 16),
    4020 => to_signed(-3811, 16),
    4021 => to_signed(-3761, 16),
    4022 => to_signed(-3711, 16),
    4023 => to_signed(-3661, 16),
    4024 => to_signed(-3611, 16),
    4025 => to_signed(-3561, 16),
    4026 => to_signed(-3511, 16),
    4027 => to_signed(-3461, 16),
    4028 => to_signed(-3411, 16),
    4029 => to_signed(-3361, 16),
    4030 => to_signed(-3311, 16),
    4031 => to_signed(-3261, 16),
    4032 => to_signed(-3211, 16),
    4033 => to_signed(-3161, 16),
    4034 => to_signed(-3111, 16),
    4035 => to_signed(-3061, 16),
    4036 => to_signed(-3011, 16),
    4037 => to_signed(-2961, 16),
    4038 => to_signed(-2911, 16),
    4039 => to_signed(-2861, 16),
    4040 => to_signed(-2811, 16),
    4041 => to_signed(-2761, 16),
    4042 => to_signed(-2711, 16),
    4043 => to_signed(-2661, 16),
    4044 => to_signed(-2610, 16),
    4045 => to_signed(-2560, 16),
    4046 => to_signed(-2510, 16),
    4047 => to_signed(-2460, 16),
    4048 => to_signed(-2410, 16),
    4049 => to_signed(-2360, 16),
    4050 => to_signed(-2310, 16),
    4051 => to_signed(-2260, 16),
    4052 => to_signed(-2209, 16),
    4053 => to_signed(-2159, 16),
    4054 => to_signed(-2109, 16),
    4055 => to_signed(-2059, 16),
    4056 => to_signed(-2009, 16),
    4057 => to_signed(-1959, 16),
    4058 => to_signed(-1908, 16),
    4059 => to_signed(-1858, 16),
    4060 => to_signed(-1808, 16),
    4061 => to_signed(-1758, 16),
    4062 => to_signed(-1708, 16),
    4063 => to_signed(-1658, 16),
    4064 => to_signed(-1607, 16),
    4065 => to_signed(-1557, 16),
    4066 => to_signed(-1507, 16),
    4067 => to_signed(-1457, 16),
    4068 => to_signed(-1406, 16),
    4069 => to_signed(-1356, 16),
    4070 => to_signed(-1306, 16),
    4071 => to_signed(-1256, 16),
    4072 => to_signed(-1206, 16),
    4073 => to_signed(-1155, 16),
    4074 => to_signed(-1105, 16),
    4075 => to_signed(-1055, 16),
    4076 => to_signed(-1005, 16),
    4077 => to_signed(-954, 16),
    4078 => to_signed(-904, 16),
    4079 => to_signed(-854, 16),
    4080 => to_signed(-804, 16),
    4081 => to_signed(-753, 16),
    4082 => to_signed(-703, 16),
    4083 => to_signed(-653, 16),
    4084 => to_signed(-603, 16),
    4085 => to_signed(-552, 16),
    4086 => to_signed(-502, 16),
    4087 => to_signed(-452, 16),
    4088 => to_signed(-402, 16),
    4089 => to_signed(-351, 16),
    4090 => to_signed(-301, 16),
    4091 => to_signed(-251, 16),
    4092 => to_signed(-201, 16),
    4093 => to_signed(-150, 16),
    4094 => to_signed(-100, 16),
    4095 => to_signed(-50, 16)
  );
end package sine_lut_pkg;
